-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(4 downto 0);
    zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_26_start: Boolean;
  signal sendOutput_CP_26_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_50_load_0_ack_1 : boolean;
  signal ptr_deref_38_load_0_req_0 : boolean;
  signal ptr_deref_38_load_0_ack_0 : boolean;
  signal ptr_deref_38_load_0_req_1 : boolean;
  signal ptr_deref_38_load_0_ack_1 : boolean;
  signal ptr_deref_50_load_0_req_0 : boolean;
  signal ptr_deref_50_load_0_ack_0 : boolean;
  signal ptr_deref_50_load_0_req_1 : boolean;
  signal type_cast_164_inst_req_0 : boolean;
  signal type_cast_164_inst_ack_0 : boolean;
  signal type_cast_164_inst_req_1 : boolean;
  signal type_cast_164_inst_ack_1 : boolean;
  signal ptr_deref_62_load_0_req_0 : boolean;
  signal ptr_deref_62_load_0_ack_0 : boolean;
  signal ptr_deref_62_load_0_req_1 : boolean;
  signal ptr_deref_62_load_0_ack_1 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal type_cast_76_inst_req_1 : boolean;
  signal type_cast_76_inst_ack_1 : boolean;
  signal if_stmt_91_branch_req_0 : boolean;
  signal if_stmt_91_branch_ack_1 : boolean;
  signal if_stmt_91_branch_ack_0 : boolean;
  signal type_cast_110_inst_req_0 : boolean;
  signal type_cast_110_inst_ack_0 : boolean;
  signal type_cast_110_inst_req_1 : boolean;
  signal type_cast_110_inst_ack_1 : boolean;
  signal array_obj_ref_145_index_offset_req_0 : boolean;
  signal array_obj_ref_145_index_offset_ack_0 : boolean;
  signal array_obj_ref_145_index_offset_req_1 : boolean;
  signal array_obj_ref_145_index_offset_ack_1 : boolean;
  signal addr_of_146_final_reg_req_0 : boolean;
  signal addr_of_146_final_reg_ack_0 : boolean;
  signal addr_of_146_final_reg_req_1 : boolean;
  signal addr_of_146_final_reg_ack_1 : boolean;
  signal ptr_deref_150_load_0_req_0 : boolean;
  signal ptr_deref_150_load_0_ack_0 : boolean;
  signal ptr_deref_150_load_0_req_1 : boolean;
  signal ptr_deref_150_load_0_ack_1 : boolean;
  signal type_cast_154_inst_req_0 : boolean;
  signal type_cast_154_inst_ack_0 : boolean;
  signal type_cast_154_inst_req_1 : boolean;
  signal type_cast_154_inst_ack_1 : boolean;
  signal type_cast_174_inst_req_0 : boolean;
  signal type_cast_174_inst_ack_0 : boolean;
  signal type_cast_174_inst_req_1 : boolean;
  signal type_cast_174_inst_ack_1 : boolean;
  signal type_cast_184_inst_req_0 : boolean;
  signal type_cast_184_inst_ack_0 : boolean;
  signal type_cast_184_inst_req_1 : boolean;
  signal type_cast_184_inst_ack_1 : boolean;
  signal type_cast_194_inst_req_0 : boolean;
  signal type_cast_194_inst_ack_0 : boolean;
  signal type_cast_194_inst_req_1 : boolean;
  signal type_cast_194_inst_ack_1 : boolean;
  signal type_cast_204_inst_req_0 : boolean;
  signal type_cast_204_inst_ack_0 : boolean;
  signal type_cast_204_inst_req_1 : boolean;
  signal type_cast_204_inst_ack_1 : boolean;
  signal type_cast_214_inst_req_0 : boolean;
  signal type_cast_214_inst_ack_0 : boolean;
  signal type_cast_214_inst_req_1 : boolean;
  signal type_cast_214_inst_ack_1 : boolean;
  signal type_cast_224_inst_req_0 : boolean;
  signal type_cast_224_inst_ack_0 : boolean;
  signal type_cast_224_inst_req_1 : boolean;
  signal type_cast_224_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_226_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_226_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_226_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_226_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_229_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_229_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_229_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_229_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_232_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_232_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_232_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_232_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_235_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_235_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_235_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_235_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_238_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_238_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_238_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_238_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_241_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_241_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_241_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_241_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_244_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_244_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_244_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_244_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_247_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_247_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_247_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_247_inst_ack_1 : boolean;
  signal if_stmt_261_branch_req_0 : boolean;
  signal if_stmt_261_branch_ack_1 : boolean;
  signal if_stmt_261_branch_ack_0 : boolean;
  signal phi_stmt_133_req_0 : boolean;
  signal type_cast_139_inst_req_0 : boolean;
  signal type_cast_139_inst_ack_0 : boolean;
  signal type_cast_139_inst_req_1 : boolean;
  signal type_cast_139_inst_ack_1 : boolean;
  signal phi_stmt_133_req_1 : boolean;
  signal phi_stmt_133_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_26_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_26: Block -- control-path 
    signal sendOutput_CP_26_elements: BooleanArray(68 downto 0);
    -- 
  begin -- 
    sendOutput_CP_26_elements(0) <= sendOutput_CP_26_start;
    sendOutput_CP_26_symbol <= sendOutput_CP_26_elements(68);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (86) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_27/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/branch_block_stmt_27__entry__
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90__entry__
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_update_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_update_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_update_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_update_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Update/cr
      -- 
    rr_89_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_89_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_38_load_0_req_0); -- 
    cr_100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_38_load_0_req_1); -- 
    rr_139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_50_load_0_req_0); -- 
    cr_150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_50_load_0_req_1); -- 
    rr_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_62_load_0_req_0); -- 
    cr_200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_62_load_0_req_1); -- 
    cr_219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => type_cast_76_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/word_access_start/word_0/ra
      -- 
    ra_90_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_38_load_0_ack_0, ack => sendOutput_CP_26_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/ptr_deref_38_Merge/$entry
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/ptr_deref_38_Merge/$exit
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/ptr_deref_38_Merge/merge_req
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/ptr_deref_38_Merge/merge_ack
      -- 
    ca_101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_38_load_0_ack_1, ack => sendOutput_CP_26_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/word_access_start/word_0/ra
      -- 
    ra_140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_50_load_0_ack_0, ack => sendOutput_CP_26_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/ptr_deref_50_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/ptr_deref_50_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/ptr_deref_50_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/ptr_deref_50_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/word_access_complete/word_0/$exit
      -- 
    ca_151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_50_load_0_ack_1, ack => sendOutput_CP_26_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/word_access_start/word_0/ra
      -- 
    ra_190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_62_load_0_ack_0, ack => sendOutput_CP_26_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/ptr_deref_62_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/ptr_deref_62_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/ptr_deref_62_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/ptr_deref_62_Merge/merge_ack
      -- 
    ca_201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_62_load_0_ack_1, ack => sendOutput_CP_26_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Sample/rr
      -- 
    rr_214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(7), ack => type_cast_76_inst_req_0); -- 
    sendOutput_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "sendOutput_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(4) & sendOutput_CP_26_elements(6) & sendOutput_CP_26_elements(2);
      gj_sendOutput_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Sample/ra
      -- 
    ra_215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_0, ack => sendOutput_CP_26_elements(8)); -- 
    -- CP-element group 9:  branch  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (13) 
      -- CP-element group 9: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90__exit__
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91__entry__
      -- CP-element group 9: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/$exit
      -- CP-element group 9: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91_dead_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91_eval_test/$entry
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91_eval_test/$exit
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91_eval_test/branch_req
      -- CP-element group 9: 	 branch_block_stmt_27/R_cmp77_92_place
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91_if_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91_else_link/$entry
      -- 
    ca_220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_1, ack => sendOutput_CP_26_elements(9)); -- 
    branch_req_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(9), ack => if_stmt_91_branch_req_0); -- 
    -- CP-element group 10:  transition  place  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	68 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 branch_block_stmt_27/if_stmt_91_if_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_27/if_stmt_91_if_link/if_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_27/entry_forx_xend
      -- CP-element group 10: 	 branch_block_stmt_27/entry_forx_xend_PhiReq/$entry
      -- CP-element group 10: 	 branch_block_stmt_27/entry_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_91_branch_ack_1, ack => sendOutput_CP_26_elements(10)); -- 
    -- CP-element group 11:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (18) 
      -- CP-element group 11: 	 branch_block_stmt_27/merge_stmt_97__exit__
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130__entry__
      -- CP-element group 11: 	 branch_block_stmt_27/if_stmt_91_else_link/$exit
      -- CP-element group 11: 	 branch_block_stmt_27/if_stmt_91_else_link/else_choice_transition
      -- CP-element group 11: 	 branch_block_stmt_27/entry_bbx_xnph
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/$entry
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_update_start_
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_27/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 11: 	 branch_block_stmt_27/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 11: 	 branch_block_stmt_27/merge_stmt_97_PhiReqMerge
      -- CP-element group 11: 	 branch_block_stmt_27/merge_stmt_97_PhiAck/$entry
      -- CP-element group 11: 	 branch_block_stmt_27/merge_stmt_97_PhiAck/$exit
      -- CP-element group 11: 	 branch_block_stmt_27/merge_stmt_97_PhiAck/dummy
      -- 
    else_choice_transition_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_91_branch_ack_0, ack => sendOutput_CP_26_elements(11)); -- 
    rr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(11), ack => type_cast_110_inst_req_0); -- 
    cr_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(11), ack => type_cast_110_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Sample/ra
      -- 
    ra_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_110_inst_ack_0, ack => sendOutput_CP_26_elements(12)); -- 
    -- CP-element group 13:  transition  place  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	62 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130__exit__
      -- CP-element group 13: 	 branch_block_stmt_27/bbx_xnph_forx_xbody
      -- CP-element group 13: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/$exit
      -- CP-element group 13: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 13: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/phi_stmt_133/$entry
      -- CP-element group 13: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/$entry
      -- 
    ca_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_110_inst_ack_1, ack => sendOutput_CP_26_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	67 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	59 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_sample_complete
      -- CP-element group 14: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Sample/ack
      -- 
    ack_285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_145_index_offset_ack_0, ack => sendOutput_CP_26_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	67 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (11) 
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_offset_calculated
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Update/ack
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_request/$entry
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_request/req
      -- 
    ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_145_index_offset_ack_1, ack => sendOutput_CP_26_elements(15)); -- 
    req_299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(15), ack => addr_of_146_final_reg_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_request/$exit
      -- CP-element group 16: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_request/ack
      -- 
    ack_300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_146_final_reg_ack_0, ack => sendOutput_CP_26_elements(16)); -- 
    -- CP-element group 17:  join  fork  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	67 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (24) 
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_complete/ack
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_word_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_root_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_address_resized
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_addr_resize/$entry
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_addr_resize/$exit
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_addr_resize/base_resize_req
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_addr_resize/base_resize_ack
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_plus_offset/$entry
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_plus_offset/$exit
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_plus_offset/sum_rename_req
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_plus_offset/sum_rename_ack
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_word_addrgen/$entry
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_word_addrgen/$exit
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_word_addrgen/root_register_req
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_word_addrgen/root_register_ack
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/word_access_start/$entry
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/word_access_start/word_0/$entry
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/word_access_start/word_0/rr
      -- 
    ack_305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_146_final_reg_ack_1, ack => sendOutput_CP_26_elements(17)); -- 
    rr_338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(17), ack => ptr_deref_150_load_0_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (5) 
      -- CP-element group 18: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/word_access_start/$exit
      -- CP-element group 18: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/word_access_start/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/word_access_start/word_0/ra
      -- 
    ra_339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_150_load_0_ack_0, ack => sendOutput_CP_26_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	67 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	24 
    -- CP-element group 19: 	26 
    -- CP-element group 19: 	28 
    -- CP-element group 19: 	30 
    -- CP-element group 19: 	32 
    -- CP-element group 19: 	34 
    -- CP-element group 19:  members (33) 
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/word_access_complete/$exit
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/word_access_complete/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/word_access_complete/word_0/ca
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/ptr_deref_150_Merge/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/ptr_deref_150_Merge/$exit
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/ptr_deref_150_Merge/merge_req
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/ptr_deref_150_Merge/merge_ack
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Sample/rr
      -- 
    ca_350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_150_load_0_ack_1, ack => sendOutput_CP_26_elements(19)); -- 
    rr_363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_154_inst_req_0); -- 
    rr_377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_164_inst_req_0); -- 
    rr_391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_174_inst_req_0); -- 
    rr_405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_184_inst_req_0); -- 
    rr_419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_194_inst_req_0); -- 
    rr_433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_204_inst_req_0); -- 
    rr_447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_214_inst_req_0); -- 
    rr_461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_224_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Sample/ra
      -- 
    ra_364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_154_inst_ack_0, ack => sendOutput_CP_26_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	67 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	56 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Update/ca
      -- 
    ca_369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_154_inst_ack_1, ack => sendOutput_CP_26_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Sample/ra
      -- 
    ra_378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_0, ack => sendOutput_CP_26_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	67 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	53 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Update/ca
      -- 
    ca_383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_1, ack => sendOutput_CP_26_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	19 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Sample/ra
      -- 
    ra_392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_174_inst_ack_0, ack => sendOutput_CP_26_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	67 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	50 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Update/ca
      -- 
    ca_397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_174_inst_ack_1, ack => sendOutput_CP_26_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	19 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Sample/ra
      -- 
    ra_406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_184_inst_ack_0, ack => sendOutput_CP_26_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	67 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	47 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Update/ca
      -- 
    ca_411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_184_inst_ack_1, ack => sendOutput_CP_26_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	19 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Sample/ra
      -- 
    ra_420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_0, ack => sendOutput_CP_26_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	67 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	44 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Update/ca
      -- 
    ca_425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_1, ack => sendOutput_CP_26_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	19 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Sample/ra
      -- 
    ra_434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_204_inst_ack_0, ack => sendOutput_CP_26_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	67 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	41 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Update/ca
      -- 
    ca_439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_204_inst_ack_1, ack => sendOutput_CP_26_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	19 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Sample/ra
      -- 
    ra_448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_0, ack => sendOutput_CP_26_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	67 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	38 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Update/ca
      -- 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_1, ack => sendOutput_CP_26_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	19 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Sample/ra
      -- 
    ra_462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_224_inst_ack_0, ack => sendOutput_CP_26_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	67 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (6) 
      -- CP-element group 35: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Sample/req
      -- 
    ca_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_224_inst_ack_1, ack => sendOutput_CP_26_elements(35)); -- 
    req_475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(35), ack => WPIPE_zeropad_output_pipe_226_inst_req_0); -- 
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_update_start_
      -- CP-element group 36: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Update/req
      -- 
    ack_476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_226_inst_ack_0, ack => sendOutput_CP_26_elements(36)); -- 
    req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(36), ack => WPIPE_zeropad_output_pipe_226_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Update/ack
      -- 
    ack_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_226_inst_ack_1, ack => sendOutput_CP_26_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	33 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Sample/req
      -- 
    req_489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(38), ack => WPIPE_zeropad_output_pipe_229_inst_req_0); -- 
    sendOutput_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(33) & sendOutput_CP_26_elements(37);
      gj_sendOutput_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_update_start_
      -- CP-element group 39: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Update/req
      -- 
    ack_490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_229_inst_ack_0, ack => sendOutput_CP_26_elements(39)); -- 
    req_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(39), ack => WPIPE_zeropad_output_pipe_229_inst_req_1); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Update/ack
      -- 
    ack_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_229_inst_ack_1, ack => sendOutput_CP_26_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	31 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Sample/req
      -- 
    req_503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(41), ack => WPIPE_zeropad_output_pipe_232_inst_req_0); -- 
    sendOutput_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(31) & sendOutput_CP_26_elements(40);
      gj_sendOutput_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_update_start_
      -- CP-element group 42: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Update/req
      -- 
    ack_504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_232_inst_ack_0, ack => sendOutput_CP_26_elements(42)); -- 
    req_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(42), ack => WPIPE_zeropad_output_pipe_232_inst_req_1); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Update/ack
      -- 
    ack_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_232_inst_ack_1, ack => sendOutput_CP_26_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	29 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Sample/req
      -- 
    req_517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(44), ack => WPIPE_zeropad_output_pipe_235_inst_req_0); -- 
    sendOutput_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(29) & sendOutput_CP_26_elements(43);
      gj_sendOutput_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_update_start_
      -- CP-element group 45: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Update/req
      -- 
    ack_518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_235_inst_ack_0, ack => sendOutput_CP_26_elements(45)); -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(45), ack => WPIPE_zeropad_output_pipe_235_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Update/ack
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_235_inst_ack_1, ack => sendOutput_CP_26_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	27 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Sample/req
      -- 
    req_531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(47), ack => WPIPE_zeropad_output_pipe_238_inst_req_0); -- 
    sendOutput_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(27) & sendOutput_CP_26_elements(46);
      gj_sendOutput_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_update_start_
      -- CP-element group 48: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Update/req
      -- 
    ack_532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_238_inst_ack_0, ack => sendOutput_CP_26_elements(48)); -- 
    req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(48), ack => WPIPE_zeropad_output_pipe_238_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Update/ack
      -- 
    ack_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_238_inst_ack_1, ack => sendOutput_CP_26_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	25 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Sample/req
      -- 
    req_545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(50), ack => WPIPE_zeropad_output_pipe_241_inst_req_0); -- 
    sendOutput_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(25) & sendOutput_CP_26_elements(49);
      gj_sendOutput_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_update_start_
      -- CP-element group 51: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Sample/ack
      -- CP-element group 51: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Update/req
      -- 
    ack_546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_241_inst_ack_0, ack => sendOutput_CP_26_elements(51)); -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(51), ack => WPIPE_zeropad_output_pipe_241_inst_req_1); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Update/ack
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_241_inst_ack_1, ack => sendOutput_CP_26_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	23 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Sample/req
      -- 
    req_559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(53), ack => WPIPE_zeropad_output_pipe_244_inst_req_0); -- 
    sendOutput_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(23) & sendOutput_CP_26_elements(52);
      gj_sendOutput_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_update_start_
      -- CP-element group 54: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Update/req
      -- 
    ack_560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_244_inst_ack_0, ack => sendOutput_CP_26_elements(54)); -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(54), ack => WPIPE_zeropad_output_pipe_244_inst_req_1); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Update/ack
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_244_inst_ack_1, ack => sendOutput_CP_26_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	21 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Sample/req
      -- 
    req_573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(56), ack => WPIPE_zeropad_output_pipe_247_inst_req_0); -- 
    sendOutput_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(21) & sendOutput_CP_26_elements(55);
      gj_sendOutput_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_update_start_
      -- CP-element group 57: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Update/req
      -- 
    ack_574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_247_inst_ack_0, ack => sendOutput_CP_26_elements(57)); -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(57), ack => WPIPE_zeropad_output_pipe_247_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Update/ack
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_247_inst_ack_1, ack => sendOutput_CP_26_elements(58)); -- 
    -- CP-element group 59:  branch  join  transition  place  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	14 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (10) 
      -- CP-element group 59: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260__exit__
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261__entry__
      -- CP-element group 59: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/$exit
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261_dead_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261_eval_test/$entry
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261_eval_test/$exit
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261_eval_test/branch_req
      -- CP-element group 59: 	 branch_block_stmt_27/R_exitcond9_262_place
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261_if_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261_else_link/$entry
      -- 
    branch_req_587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(59), ack => if_stmt_261_branch_req_0); -- 
    sendOutput_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(14) & sendOutput_CP_26_elements(58);
      gj_sendOutput_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  merge  transition  place  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	68 
    -- CP-element group 60:  members (13) 
      -- CP-element group 60: 	 branch_block_stmt_27/merge_stmt_267__exit__
      -- CP-element group 60: 	 branch_block_stmt_27/forx_xendx_xloopexit_forx_xend
      -- CP-element group 60: 	 branch_block_stmt_27/if_stmt_261_if_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_27/if_stmt_261_if_link/if_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_27/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 60: 	 branch_block_stmt_27/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_27/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_27/merge_stmt_267_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_27/merge_stmt_267_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_27/merge_stmt_267_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_27/merge_stmt_267_PhiAck/dummy
      -- CP-element group 60: 	 branch_block_stmt_27/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_27/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_261_branch_ack_1, ack => sendOutput_CP_26_elements(60)); -- 
    -- CP-element group 61:  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: 	64 
    -- CP-element group 61:  members (12) 
      -- CP-element group 61: 	 branch_block_stmt_27/if_stmt_261_else_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_27/if_stmt_261_else_link/else_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Update/cr
      -- 
    else_choice_transition_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_261_branch_ack_0, ack => sendOutput_CP_26_elements(61)); -- 
    rr_640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(61), ack => type_cast_139_inst_req_0); -- 
    cr_645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(61), ack => type_cast_139_inst_req_1); -- 
    -- CP-element group 62:  transition  output  delay-element  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	13 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	66 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/phi_stmt_133/$exit
      -- CP-element group 62: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/$exit
      -- CP-element group 62: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_137_konst_delay_trans
      -- CP-element group 62: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_req
      -- 
    phi_stmt_133_req_621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_133_req_621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(62), ack => phi_stmt_133_req_0); -- 
    -- Element group sendOutput_CP_26_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => sendOutput_CP_26_elements(13), ack => sendOutput_CP_26_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Sample/ra
      -- 
    ra_641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_0, ack => sendOutput_CP_26_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	61 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Update/ca
      -- 
    ca_646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_1, ack => sendOutput_CP_26_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/$exit
      -- CP-element group 65: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/$exit
      -- CP-element group 65: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/$exit
      -- CP-element group 65: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/$exit
      -- CP-element group 65: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_req
      -- 
    phi_stmt_133_req_647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_133_req_647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(65), ack => phi_stmt_133_req_1); -- 
    sendOutput_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(63) & sendOutput_CP_26_elements(64);
      gj_sendOutput_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  merge  transition  place  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	62 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_27/merge_stmt_132_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_27/merge_stmt_132_PhiAck/$entry
      -- 
    sendOutput_CP_26_elements(66) <= OrReduce(sendOutput_CP_26_elements(62) & sendOutput_CP_26_elements(65));
    -- CP-element group 67:  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	14 
    -- CP-element group 67: 	15 
    -- CP-element group 67: 	17 
    -- CP-element group 67: 	19 
    -- CP-element group 67: 	21 
    -- CP-element group 67: 	23 
    -- CP-element group 67: 	25 
    -- CP-element group 67: 	27 
    -- CP-element group 67: 	29 
    -- CP-element group 67: 	31 
    -- CP-element group 67: 	33 
    -- CP-element group 67: 	35 
    -- CP-element group 67:  members (53) 
      -- CP-element group 67: 	 branch_block_stmt_27/merge_stmt_132__exit__
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260__entry__
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_resized_1
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_scaled_1
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_computed_1
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_resize_1/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_resize_1/$exit
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_resize_1/index_resize_req
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_resize_1/index_resize_ack
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_scale_1/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_scale_1/$exit
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_scale_1/scale_rename_req
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_scale_1/scale_rename_ack
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_update_start
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Sample/req
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Update/req
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_complete/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_complete/req
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/word_access_complete/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/word_access_complete/word_0/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/word_access_complete/word_0/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/merge_stmt_132_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_27/merge_stmt_132_PhiAck/phi_stmt_133_ack
      -- 
    phi_stmt_133_ack_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_133_ack_0, ack => sendOutput_CP_26_elements(67)); -- 
    cr_382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_164_inst_req_1); -- 
    req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => array_obj_ref_145_index_offset_req_0); -- 
    req_289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => array_obj_ref_145_index_offset_req_1); -- 
    req_304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => addr_of_146_final_reg_req_1); -- 
    cr_349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => ptr_deref_150_load_0_req_1); -- 
    cr_368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_154_inst_req_1); -- 
    cr_396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_174_inst_req_1); -- 
    cr_410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_184_inst_req_1); -- 
    cr_424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_194_inst_req_1); -- 
    cr_438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_204_inst_req_1); -- 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_214_inst_req_1); -- 
    cr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_224_inst_req_1); -- 
    -- CP-element group 68:  merge  transition  place  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	10 
    -- CP-element group 68: 	60 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 $exit
      -- CP-element group 68: 	 branch_block_stmt_27/$exit
      -- CP-element group 68: 	 branch_block_stmt_27/branch_block_stmt_27__exit__
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_269__exit__
      -- CP-element group 68: 	 branch_block_stmt_27/return__
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_271__exit__
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_269_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_269_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_269_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_269_PhiAck/dummy
      -- CP-element group 68: 	 branch_block_stmt_27/return___PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_27/return___PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_271_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_271_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_271_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_271_PhiAck/dummy
      -- 
    sendOutput_CP_26_elements(68) <= OrReduce(sendOutput_CP_26_elements(10) & sendOutput_CP_26_elements(60));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_144_resized : std_logic_vector(13 downto 0);
    signal R_indvar_144_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_145_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_145_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_145_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_145_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_145_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_145_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_147 : std_logic_vector(31 downto 0);
    signal cmp77_90 : std_logic_vector(0 downto 0);
    signal conv14_155 : std_logic_vector(7 downto 0);
    signal conv20_165 : std_logic_vector(7 downto 0);
    signal conv26_175 : std_logic_vector(7 downto 0);
    signal conv32_185 : std_logic_vector(7 downto 0);
    signal conv38_195 : std_logic_vector(7 downto 0);
    signal conv44_205 : std_logic_vector(7 downto 0);
    signal conv50_215 : std_logic_vector(7 downto 0);
    signal conv56_225 : std_logic_vector(7 downto 0);
    signal conv_77 : std_logic_vector(63 downto 0);
    signal exitcond9_260 : std_logic_vector(0 downto 0);
    signal iNsTr_0_35 : std_logic_vector(31 downto 0);
    signal iNsTr_1_47 : std_logic_vector(31 downto 0);
    signal iNsTr_2_59 : std_logic_vector(31 downto 0);
    signal indvar_133 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_255 : std_logic_vector(63 downto 0);
    signal mul3_73 : std_logic_vector(31 downto 0);
    signal mul_68 : std_logic_vector(31 downto 0);
    signal ptr_deref_150_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_150_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_150_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_150_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_150_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_38_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_38_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_38_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_38_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_38_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_50_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_50_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_50_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_50_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_50_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_62_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_62_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_62_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_62_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_62_word_offset_0 : std_logic_vector(6 downto 0);
    signal shr17_161 : std_logic_vector(63 downto 0);
    signal shr23_171 : std_logic_vector(63 downto 0);
    signal shr29_181 : std_logic_vector(63 downto 0);
    signal shr35_191 : std_logic_vector(63 downto 0);
    signal shr41_201 : std_logic_vector(63 downto 0);
    signal shr47_211 : std_logic_vector(63 downto 0);
    signal shr53_221 : std_logic_vector(63 downto 0);
    signal shr76x_xmask_83 : std_logic_vector(63 downto 0);
    signal tmp11_151 : std_logic_vector(63 downto 0);
    signal tmp1_51 : std_logic_vector(31 downto 0);
    signal tmp2_63 : std_logic_vector(31 downto 0);
    signal tmp3_102 : std_logic_vector(31 downto 0);
    signal tmp4_107 : std_logic_vector(31 downto 0);
    signal tmp5_111 : std_logic_vector(63 downto 0);
    signal tmp6_117 : std_logic_vector(63 downto 0);
    signal tmp7_123 : std_logic_vector(0 downto 0);
    signal tmp_39 : std_logic_vector(31 downto 0);
    signal type_cast_115_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_121_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_128_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_137_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_139_wire : std_logic_vector(63 downto 0);
    signal type_cast_159_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_169_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_179_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_189_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_199_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_209_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_219_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_253_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_81_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_87_wire_constant : std_logic_vector(63 downto 0);
    signal umax8_130 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_145_constant_part_of_offset <= "00000000000000";
    array_obj_ref_145_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_145_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_145_resized_base_address <= "00000000000000";
    iNsTr_0_35 <= "00000000000000000000000000000011";
    iNsTr_1_47 <= "00000000000000000000000000000100";
    iNsTr_2_59 <= "00000000000000000000000000000101";
    ptr_deref_150_word_offset_0 <= "00000000000000";
    ptr_deref_38_word_offset_0 <= "0000000";
    ptr_deref_50_word_offset_0 <= "0000000";
    ptr_deref_62_word_offset_0 <= "0000000";
    type_cast_115_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_121_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_128_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_137_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_159_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_169_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_179_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_189_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_199_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_209_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_219_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_253_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_81_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_87_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_133: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_137_wire_constant & type_cast_139_wire;
      req <= phi_stmt_133_req_0 & phi_stmt_133_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_133",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_133_ack_0,
          idata => idata,
          odata => indvar_133,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_133
    -- flow-through select operator MUX_129_inst
    umax8_130 <= tmp6_117 when (tmp7_123(0) /=  '0') else type_cast_128_wire_constant;
    addr_of_146_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_146_final_reg_req_0;
      addr_of_146_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_146_final_reg_req_1;
      addr_of_146_final_reg_ack_1<= rack(0);
      addr_of_146_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_146_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_145_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_147,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_110_inst_req_0;
      type_cast_110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_110_inst_req_1;
      type_cast_110_inst_ack_1<= rack(0);
      type_cast_110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp5_111,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_139_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_139_inst_req_0;
      type_cast_139_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_139_inst_req_1;
      type_cast_139_inst_ack_1<= rack(0);
      type_cast_139_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_139_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_255,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_139_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_154_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_154_inst_req_0;
      type_cast_154_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_154_inst_req_1;
      type_cast_154_inst_ack_1<= rack(0);
      type_cast_154_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_154_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp11_151,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv14_155,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_164_inst_req_0;
      type_cast_164_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_164_inst_req_1;
      type_cast_164_inst_ack_1<= rack(0);
      type_cast_164_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_164_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr17_161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_174_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_174_inst_req_0;
      type_cast_174_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_174_inst_req_1;
      type_cast_174_inst_ack_1<= rack(0);
      type_cast_174_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_174_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr23_171,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_175,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_184_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_184_inst_req_0;
      type_cast_184_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_184_inst_req_1;
      type_cast_184_inst_ack_1<= rack(0);
      type_cast_184_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_184_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr29_181,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_185,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_194_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_194_inst_req_0;
      type_cast_194_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_194_inst_req_1;
      type_cast_194_inst_ack_1<= rack(0);
      type_cast_194_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_194_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr35_191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_195,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_204_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_204_inst_req_0;
      type_cast_204_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_204_inst_req_1;
      type_cast_204_inst_ack_1<= rack(0);
      type_cast_204_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_204_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr41_201,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_205,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_214_inst_req_0;
      type_cast_214_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_214_inst_req_1;
      type_cast_214_inst_ack_1<= rack(0);
      type_cast_214_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_214_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr47_211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_215,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_224_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_224_inst_req_0;
      type_cast_224_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_224_inst_req_1;
      type_cast_224_inst_ack_1<= rack(0);
      type_cast_224_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_224_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr53_221,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_225,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_76_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_76_inst_req_0;
      type_cast_76_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_76_inst_req_1;
      type_cast_76_inst_ack_1<= rack(0);
      type_cast_76_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_76_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul3_73,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_77,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_145_index_1_rename
    process(R_indvar_144_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_144_resized;
      ov(13 downto 0) := iv;
      R_indvar_144_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_145_index_1_resize
    process(indvar_133) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_133;
      ov := iv(13 downto 0);
      R_indvar_144_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_145_root_address_inst
    process(array_obj_ref_145_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_145_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_145_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_150_addr_0
    process(ptr_deref_150_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_150_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_150_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_150_base_resize
    process(arrayidx_147) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_147;
      ov := iv(13 downto 0);
      ptr_deref_150_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_150_gather_scatter
    process(ptr_deref_150_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_150_data_0;
      ov(63 downto 0) := iv;
      tmp11_151 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_150_root_address_inst
    process(ptr_deref_150_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_150_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_150_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_38_addr_0
    process(ptr_deref_38_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_38_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_38_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_38_base_resize
    process(iNsTr_0_35) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_35;
      ov := iv(6 downto 0);
      ptr_deref_38_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_38_gather_scatter
    process(ptr_deref_38_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_38_data_0;
      ov(31 downto 0) := iv;
      tmp_39 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_38_root_address_inst
    process(ptr_deref_38_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_38_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_38_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_50_addr_0
    process(ptr_deref_50_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_50_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_50_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_50_base_resize
    process(iNsTr_1_47) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_47;
      ov := iv(6 downto 0);
      ptr_deref_50_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_50_gather_scatter
    process(ptr_deref_50_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_50_data_0;
      ov(31 downto 0) := iv;
      tmp1_51 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_50_root_address_inst
    process(ptr_deref_50_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_50_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_50_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_62_addr_0
    process(ptr_deref_62_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_62_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_62_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_62_base_resize
    process(iNsTr_2_59) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_59;
      ov := iv(6 downto 0);
      ptr_deref_62_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_62_gather_scatter
    process(ptr_deref_62_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_62_data_0;
      ov(31 downto 0) := iv;
      tmp2_63 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_62_root_address_inst
    process(ptr_deref_62_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_62_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_62_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_261_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond9_260;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_261_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_261_branch_req_0,
          ack0 => if_stmt_261_branch_ack_0,
          ack1 => if_stmt_261_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_91_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_90;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_91_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_91_branch_req_0,
          ack0 => if_stmt_91_branch_ack_0,
          ack1 => if_stmt_91_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_254_inst
    process(indvar_133) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_133, type_cast_253_wire_constant, tmp_var);
      indvarx_xnext_255 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_82_inst
    process(conv_77) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv_77, type_cast_81_wire_constant, tmp_var);
      shr76x_xmask_83 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_259_inst
    process(indvarx_xnext_255, umax8_130) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_255, umax8_130, tmp_var);
      exitcond9_260 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_88_inst
    process(shr76x_xmask_83) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr76x_xmask_83, type_cast_87_wire_constant, tmp_var);
      cmp77_90 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_116_inst
    process(tmp5_111) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_111, type_cast_115_wire_constant, tmp_var);
      tmp6_117 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_160_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_159_wire_constant, tmp_var);
      shr17_161 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_170_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_169_wire_constant, tmp_var);
      shr23_171 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_180_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_179_wire_constant, tmp_var);
      shr29_181 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_190_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_189_wire_constant, tmp_var);
      shr35_191 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_200_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_199_wire_constant, tmp_var);
      shr41_201 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_210_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_209_wire_constant, tmp_var);
      shr47_211 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_220_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_219_wire_constant, tmp_var);
      shr53_221 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_101_inst
    process(tmp1_51, tmp_39) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_51, tmp_39, tmp_var);
      tmp3_102 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_106_inst
    process(tmp3_102, tmp2_63) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp3_102, tmp2_63, tmp_var);
      tmp4_107 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_67_inst
    process(tmp1_51, tmp_39) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_51, tmp_39, tmp_var);
      mul_68 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_72_inst
    process(mul_68, tmp2_63) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_68, tmp2_63, tmp_var);
      mul3_73 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_122_inst
    process(tmp6_117) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp6_117, type_cast_121_wire_constant, tmp_var);
      tmp7_123 <= tmp_var; --
    end process;
    -- shared split operator group (17) : array_obj_ref_145_index_offset 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_144_scaled;
      array_obj_ref_145_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_145_index_offset_req_0;
      array_obj_ref_145_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_145_index_offset_req_1;
      array_obj_ref_145_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_17_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared load operator group (0) : ptr_deref_150_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_150_load_0_req_0;
      ptr_deref_150_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_150_load_0_req_1;
      ptr_deref_150_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_150_word_address_0;
      ptr_deref_150_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_38_load_0 ptr_deref_50_load_0 ptr_deref_62_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_38_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_50_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_62_load_0_req_0;
      ptr_deref_38_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_50_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_62_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_38_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_50_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_62_load_0_req_1;
      ptr_deref_38_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_50_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_62_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_38_word_address_0 & ptr_deref_50_word_address_0 & ptr_deref_62_word_address_0;
      ptr_deref_38_data_0 <= data_out(95 downto 64);
      ptr_deref_50_data_0 <= data_out(63 downto 32);
      ptr_deref_62_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(6 downto 0),
          mtag => memory_space_6_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(31 downto 0),
          mtag => memory_space_6_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared outport operator group (0) : WPIPE_zeropad_output_pipe_226_inst WPIPE_zeropad_output_pipe_229_inst WPIPE_zeropad_output_pipe_232_inst WPIPE_zeropad_output_pipe_235_inst WPIPE_zeropad_output_pipe_238_inst WPIPE_zeropad_output_pipe_241_inst WPIPE_zeropad_output_pipe_244_inst WPIPE_zeropad_output_pipe_247_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_zeropad_output_pipe_226_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_zeropad_output_pipe_229_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_zeropad_output_pipe_232_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_zeropad_output_pipe_235_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_zeropad_output_pipe_238_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_zeropad_output_pipe_241_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_zeropad_output_pipe_244_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_zeropad_output_pipe_247_inst_req_0;
      WPIPE_zeropad_output_pipe_226_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_229_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_232_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_235_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_238_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_241_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_244_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_247_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_zeropad_output_pipe_226_inst_req_1;
      update_req_unguarded(6) <= WPIPE_zeropad_output_pipe_229_inst_req_1;
      update_req_unguarded(5) <= WPIPE_zeropad_output_pipe_232_inst_req_1;
      update_req_unguarded(4) <= WPIPE_zeropad_output_pipe_235_inst_req_1;
      update_req_unguarded(3) <= WPIPE_zeropad_output_pipe_238_inst_req_1;
      update_req_unguarded(2) <= WPIPE_zeropad_output_pipe_241_inst_req_1;
      update_req_unguarded(1) <= WPIPE_zeropad_output_pipe_244_inst_req_1;
      update_req_unguarded(0) <= WPIPE_zeropad_output_pipe_247_inst_req_1;
      WPIPE_zeropad_output_pipe_226_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_229_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_232_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_235_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_238_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_241_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_244_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_247_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv56_225 & conv50_215 & conv44_205 & conv38_195 & conv32_185 & conv26_175 & conv20_165 & conv14_155;
      zeropad_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "zeropad_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      zeropad_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "zeropad_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => zeropad_output_pipe_pipe_write_req(0),
          oack => zeropad_output_pipe_pipe_write_ack(0),
          odata => zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(4 downto 0);
    zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal ret_val_x_x_update_enable: Boolean;
  signal testConfigure_CP_684_start: Boolean;
  signal testConfigure_CP_684_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal STORE_row_high_326_store_0_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_330_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_330_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_307_inst_ack_1 : boolean;
  signal type_cast_595_inst_req_1 : boolean;
  signal type_cast_595_inst_ack_0 : boolean;
  signal type_cast_595_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_609_inst_req_1 : boolean;
  signal ptr_deref_320_store_0_ack_0 : boolean;
  signal type_cast_595_inst_ack_1 : boolean;
  signal type_cast_528_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_330_inst_req_0 : boolean;
  signal type_cast_649_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_330_inst_ack_0 : boolean;
  signal type_cast_528_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_307_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_290_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_324_inst_req_0 : boolean;
  signal STORE_row_high_326_store_0_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_307_inst_ack_0 : boolean;
  signal STORE_row_high_326_store_0_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_307_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_290_inst_ack_0 : boolean;
  signal type_cast_294_inst_ack_1 : boolean;
  signal type_cast_294_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_324_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_555_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_290_inst_req_0 : boolean;
  signal type_cast_294_inst_ack_0 : boolean;
  signal type_cast_294_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_609_inst_ack_1 : boolean;
  signal type_cast_311_inst_ack_1 : boolean;
  signal type_cast_311_inst_req_1 : boolean;
  signal ptr_deref_285_store_0_ack_1 : boolean;
  signal ptr_deref_303_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_609_inst_req_0 : boolean;
  signal ptr_deref_285_store_0_req_1 : boolean;
  signal ptr_deref_303_store_0_req_1 : boolean;
  signal type_cast_613_inst_req_0 : boolean;
  signal type_cast_528_inst_req_1 : boolean;
  signal ptr_deref_320_store_0_req_0 : boolean;
  signal ptr_deref_303_store_0_ack_0 : boolean;
  signal ptr_deref_285_store_0_ack_0 : boolean;
  signal type_cast_613_inst_ack_0 : boolean;
  signal ptr_deref_285_store_0_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_609_inst_ack_0 : boolean;
  signal ptr_deref_303_store_0_req_0 : boolean;
  signal type_cast_631_inst_req_0 : boolean;
  signal type_cast_682_inst_req_0 : boolean;
  signal type_cast_682_inst_ack_1 : boolean;
  signal phi_stmt_508_req_0 : boolean;
  signal array_obj_ref_520_index_offset_req_0 : boolean;
  signal type_cast_311_inst_ack_0 : boolean;
  signal type_cast_311_inst_req_0 : boolean;
  signal ptr_deref_320_store_0_ack_1 : boolean;
  signal ptr_deref_320_store_0_req_1 : boolean;
  signal type_cast_631_inst_ack_0 : boolean;
  signal type_cast_528_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_324_inst_ack_1 : boolean;
  signal STORE_row_high_326_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_324_inst_req_1 : boolean;
  signal array_obj_ref_520_index_offset_ack_0 : boolean;
  signal type_cast_613_inst_req_1 : boolean;
  signal type_cast_613_inst_ack_1 : boolean;
  signal addr_of_521_final_reg_req_0 : boolean;
  signal addr_of_521_final_reg_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_627_inst_req_0 : boolean;
  signal type_cast_631_inst_req_1 : boolean;
  signal type_cast_631_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_537_inst_req_0 : boolean;
  signal addr_of_521_final_reg_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_537_inst_ack_0 : boolean;
  signal addr_of_521_final_reg_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_627_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_627_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_537_inst_req_1 : boolean;
  signal type_cast_514_inst_ack_1 : boolean;
  signal if_stmt_671_branch_req_0 : boolean;
  signal phi_stmt_508_req_1 : boolean;
  signal type_cast_514_inst_req_1 : boolean;
  signal type_cast_514_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_537_inst_ack_1 : boolean;
  signal type_cast_514_inst_ack_0 : boolean;
  signal array_obj_ref_520_index_offset_req_1 : boolean;
  signal array_obj_ref_520_index_offset_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_627_inst_ack_1 : boolean;
  signal type_cast_682_inst_req_1 : boolean;
  signal type_cast_541_inst_req_0 : boolean;
  signal type_cast_541_inst_ack_0 : boolean;
  signal type_cast_541_inst_req_1 : boolean;
  signal if_stmt_671_branch_ack_0 : boolean;
  signal type_cast_682_inst_ack_0 : boolean;
  signal type_cast_541_inst_ack_1 : boolean;
  signal type_cast_559_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_290_inst_ack_1 : boolean;
  signal type_cast_649_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_555_inst_req_1 : boolean;
  signal STORE_col_high_332_store_0_req_0 : boolean;
  signal STORE_col_high_332_store_0_ack_0 : boolean;
  signal STORE_col_high_332_store_0_req_1 : boolean;
  signal STORE_col_high_332_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_336_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_336_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_336_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_336_inst_ack_1 : boolean;
  signal ptr_deref_657_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_591_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_591_inst_req_1 : boolean;
  signal type_cast_649_inst_ack_0 : boolean;
  signal STORE_depth_high_338_store_0_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_591_inst_ack_0 : boolean;
  signal STORE_depth_high_338_store_0_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_555_inst_ack_0 : boolean;
  signal STORE_depth_high_338_store_0_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_591_inst_req_0 : boolean;
  signal STORE_depth_high_338_store_0_ack_1 : boolean;
  signal ptr_deref_657_store_0_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_342_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_342_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_342_inst_req_1 : boolean;
  signal type_cast_649_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_342_inst_ack_1 : boolean;
  signal if_stmt_671_branch_ack_1 : boolean;
  signal type_cast_577_inst_ack_1 : boolean;
  signal type_cast_577_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_555_inst_req_0 : boolean;
  signal STORE_pad_344_store_0_req_0 : boolean;
  signal STORE_pad_344_store_0_ack_0 : boolean;
  signal STORE_pad_344_store_0_req_1 : boolean;
  signal type_cast_577_inst_ack_0 : boolean;
  signal STORE_pad_344_store_0_ack_1 : boolean;
  signal type_cast_577_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_348_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_348_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_524_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_348_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_348_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_524_inst_req_1 : boolean;
  signal type_cast_352_inst_req_0 : boolean;
  signal type_cast_352_inst_ack_0 : boolean;
  signal type_cast_352_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_645_inst_ack_1 : boolean;
  signal type_cast_352_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_573_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_573_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_573_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_645_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_524_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_573_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_524_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_645_inst_ack_0 : boolean;
  signal ptr_deref_363_store_0_req_0 : boolean;
  signal ptr_deref_363_store_0_ack_0 : boolean;
  signal ptr_deref_363_store_0_req_1 : boolean;
  signal ptr_deref_363_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_645_inst_req_0 : boolean;
  signal type_cast_559_inst_ack_1 : boolean;
  signal type_cast_559_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_ack_1 : boolean;
  signal ptr_deref_657_store_0_ack_0 : boolean;
  signal type_cast_559_inst_ack_0 : boolean;
  signal ptr_deref_657_store_0_req_0 : boolean;
  signal type_cast_371_inst_req_0 : boolean;
  signal type_cast_371_inst_ack_0 : boolean;
  signal type_cast_371_inst_req_1 : boolean;
  signal type_cast_371_inst_ack_1 : boolean;
  signal ptr_deref_382_store_0_req_0 : boolean;
  signal ptr_deref_382_store_0_ack_0 : boolean;
  signal ptr_deref_382_store_0_req_1 : boolean;
  signal ptr_deref_382_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_386_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_386_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_386_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_386_inst_ack_1 : boolean;
  signal type_cast_390_inst_req_0 : boolean;
  signal type_cast_390_inst_ack_0 : boolean;
  signal type_cast_390_inst_req_1 : boolean;
  signal type_cast_390_inst_ack_1 : boolean;
  signal ptr_deref_401_store_0_req_0 : boolean;
  signal ptr_deref_401_store_0_ack_0 : boolean;
  signal ptr_deref_401_store_0_req_1 : boolean;
  signal ptr_deref_401_store_0_ack_1 : boolean;
  signal ptr_deref_414_load_0_req_0 : boolean;
  signal ptr_deref_414_load_0_ack_0 : boolean;
  signal ptr_deref_414_load_0_req_1 : boolean;
  signal ptr_deref_414_load_0_ack_1 : boolean;
  signal ptr_deref_426_load_0_req_0 : boolean;
  signal ptr_deref_426_load_0_ack_0 : boolean;
  signal ptr_deref_426_load_0_req_1 : boolean;
  signal ptr_deref_426_load_0_ack_1 : boolean;
  signal ptr_deref_438_load_0_req_0 : boolean;
  signal ptr_deref_438_load_0_ack_0 : boolean;
  signal ptr_deref_438_load_0_req_1 : boolean;
  signal ptr_deref_438_load_0_ack_1 : boolean;
  signal type_cast_452_inst_req_0 : boolean;
  signal type_cast_452_inst_ack_0 : boolean;
  signal type_cast_452_inst_req_1 : boolean;
  signal type_cast_452_inst_ack_1 : boolean;
  signal if_stmt_466_branch_req_0 : boolean;
  signal if_stmt_466_branch_ack_1 : boolean;
  signal if_stmt_466_branch_ack_0 : boolean;
  signal type_cast_485_inst_req_0 : boolean;
  signal type_cast_485_inst_ack_0 : boolean;
  signal type_cast_485_inst_req_1 : boolean;
  signal type_cast_485_inst_ack_1 : boolean;
  signal phi_stmt_508_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_684_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_684_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_684_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_684_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_684: Block -- control-path 
    signal testConfigure_CP_684_elements: BooleanArray(132 downto 0);
    -- 
  begin -- 
    testConfigure_CP_684_elements(0) <= testConfigure_CP_684_start;
    testConfigure_CP_684_symbol <= testConfigure_CP_684_elements(125);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	47 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	58 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	61 
    -- CP-element group 0: 	63 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	66 
    -- CP-element group 0: 	26 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	54 
    -- CP-element group 0: 	55 
    -- CP-element group 0: 	31 
    -- CP-element group 0: 	34 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	50 
    -- CP-element group 0: 	14 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	43 
    -- CP-element group 0: 	19 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0:  members (252) 
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465__entry__
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/ptr_deref_285_Split/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/branch_block_stmt_277__entry__
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/ptr_deref_285_Split/split_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/ptr_deref_285_Split/split_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/ptr_deref_285_Split/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_address_resized
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Update/cr
      -- 
    cr_968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => STORE_row_high_326_store_0_req_1); -- 
    cr_793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_294_inst_req_1); -- 
    rr_774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => RPIPE_zeropad_input_pipe_290_inst_req_0); -- 
    cr_871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_311_inst_req_1); -- 
    cr_765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_285_store_0_req_1); -- 
    cr_843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_303_store_0_req_1); -- 
    rr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_285_store_0_req_0); -- 
    cr_921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_320_store_0_req_1); -- 
    cr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => STORE_col_high_332_store_0_req_1); -- 
    cr_1062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => STORE_depth_high_338_store_0_req_1); -- 
    cr_1109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => STORE_pad_344_store_0_req_1); -- 
    cr_1137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_352_inst_req_1); -- 
    cr_1187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_363_store_0_req_1); -- 
    cr_1215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_371_inst_req_1); -- 
    cr_1265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_382_store_0_req_1); -- 
    cr_1293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_390_inst_req_1); -- 
    cr_1343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_401_store_0_req_1); -- 
    cr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_414_load_0_req_1); -- 
    cr_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_426_load_0_req_1); -- 
    cr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_438_load_0_req_1); -- 
    cr_1507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_452_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	70 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/$exit
      -- 
    ra_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_285_store_0_ack_0, ack => testConfigure_CP_684_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	77 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_update_completed_
      -- 
    ca_766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_285_store_0_ack_1, ack => testConfigure_CP_684_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_update_start_
      -- CP-element group 3: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_sample_completed_
      -- 
    ra_775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_290_inst_ack_0, ack => testConfigure_CP_684_elements(3)); -- 
    cr_779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(3), ack => RPIPE_zeropad_input_pipe_290_inst_req_1); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Update/ca
      -- 
    ca_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_290_inst_ack_1, ack => testConfigure_CP_684_elements(4)); -- 
    rr_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(4), ack => RPIPE_zeropad_input_pipe_307_inst_req_0); -- 
    rr_788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(4), ack => type_cast_294_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_sample_completed_
      -- 
    ra_789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_294_inst_ack_0, ack => testConfigure_CP_684_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_update_completed_
      -- 
    ca_794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_294_inst_ack_1, ack => testConfigure_CP_684_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	70 
    -- CP-element group 7: 	0 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/word_access_start/word_0/rr
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/word_access_start/word_0/$entry
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/word_access_start/$entry
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/ptr_deref_303_Split/split_ack
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/ptr_deref_303_Split/split_req
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/ptr_deref_303_Split/$exit
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/ptr_deref_303_Split/$entry
      -- 
    rr_832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(7), ack => ptr_deref_303_store_0_req_0); -- 
    testConfigure_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(70) & testConfigure_CP_684_elements(0) & testConfigure_CP_684_elements(6);
      gj_testConfigure_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	71 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/word_access_start/word_0/ra
      -- CP-element group 8: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/word_access_start/$exit
      -- 
    ra_833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_303_store_0_ack_0, ack => testConfigure_CP_684_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	77 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/word_access_complete/$exit
      -- CP-element group 9: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_update_completed_
      -- 
    ca_844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_303_store_0_ack_1, ack => testConfigure_CP_684_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_update_start_
      -- CP-element group 10: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_sample_completed_
      -- 
    ra_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_307_inst_ack_0, ack => testConfigure_CP_684_elements(10)); -- 
    cr_857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(10), ack => RPIPE_zeropad_input_pipe_307_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_sample_start_
      -- 
    ca_858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_307_inst_ack_1, ack => testConfigure_CP_684_elements(11)); -- 
    rr_866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(11), ack => type_cast_311_inst_req_0); -- 
    rr_930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(11), ack => RPIPE_zeropad_input_pipe_324_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_sample_completed_
      -- 
    ra_867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_311_inst_ack_0, ack => testConfigure_CP_684_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_update_completed_
      -- 
    ca_872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_311_inst_ack_1, ack => testConfigure_CP_684_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: 	71 
    -- CP-element group 14: 	0 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/word_access_start/word_0/rr
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/word_access_start/word_0/$entry
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/word_access_start/$entry
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/ptr_deref_320_Split/split_ack
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/ptr_deref_320_Split/split_req
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/ptr_deref_320_Split/$exit
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/ptr_deref_320_Split/$entry
      -- 
    rr_910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(14), ack => ptr_deref_320_store_0_req_0); -- 
    testConfigure_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(13) & testConfigure_CP_684_elements(71) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	72 
    -- CP-element group 15: 	73 
    -- CP-element group 15: 	74 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/word_access_start/word_0/ra
      -- CP-element group 15: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/$exit
      -- 
    ra_911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_320_store_0_ack_0, ack => testConfigure_CP_684_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	77 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/word_access_complete/word_0/ca
      -- 
    ca_922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_320_store_0_ack_1, ack => testConfigure_CP_684_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_update_start_
      -- CP-element group 17: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Update/cr
      -- 
    ra_931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_324_inst_ack_0, ack => testConfigure_CP_684_elements(17)); -- 
    cr_935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(17), ack => RPIPE_zeropad_input_pipe_324_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	22 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Update/ca
      -- 
    ca_936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_324_inst_ack_1, ack => testConfigure_CP_684_elements(18)); -- 
    rr_977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(18), ack => RPIPE_zeropad_input_pipe_330_inst_req_0); -- 
    -- CP-element group 19:  join  transition  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	0 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/word_access_start/word_0/rr
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/word_access_start/word_0/$entry
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/word_access_start/$entry
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/STORE_row_high_326_Split/split_ack
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/STORE_row_high_326_Split/split_req
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/STORE_row_high_326_Split/$exit
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/STORE_row_high_326_Split/$entry
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/$entry
      -- 
    rr_957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(19), ack => STORE_row_high_326_store_0_req_0); -- 
    testConfigure_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(0) & testConfigure_CP_684_elements(18);
      gj_testConfigure_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/word_access_start/word_0/ra
      -- CP-element group 20: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/word_access_start/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/word_access_start/$exit
      -- CP-element group 20: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/$exit
      -- 
    ra_958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_row_high_326_store_0_ack_0, ack => testConfigure_CP_684_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	77 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/word_access_complete/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/word_access_complete/$exit
      -- CP-element group 21: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/word_access_complete/word_0/ca
      -- 
    ca_969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_row_high_326_store_0_ack_1, ack => testConfigure_CP_684_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	18 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_update_start_
      -- CP-element group 22: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Sample/ra
      -- 
    ra_978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_330_inst_ack_0, ack => testConfigure_CP_684_elements(22)); -- 
    cr_982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(22), ack => RPIPE_zeropad_input_pipe_330_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	27 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Sample/rr
      -- 
    ca_983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_330_inst_ack_1, ack => testConfigure_CP_684_elements(23)); -- 
    rr_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(23), ack => RPIPE_zeropad_input_pipe_336_inst_req_0); -- 
    -- CP-element group 24:  join  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/STORE_col_high_332_Split/$entry
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/STORE_col_high_332_Split/$exit
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/STORE_col_high_332_Split/split_req
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/STORE_col_high_332_Split/split_ack
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/word_access_start/$entry
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/word_access_start/word_0/$entry
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/word_access_start/word_0/rr
      -- 
    rr_1004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(24), ack => STORE_col_high_332_store_0_req_0); -- 
    testConfigure_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(23) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/word_access_start/word_0/ra
      -- 
    ra_1005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_col_high_332_store_0_ack_0, ack => testConfigure_CP_684_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	0 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	77 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/word_access_complete/word_0/ca
      -- 
    ca_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_col_high_332_store_0_ack_1, ack => testConfigure_CP_684_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	23 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_update_start_
      -- CP-element group 27: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Update/cr
      -- 
    ra_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_336_inst_ack_0, ack => testConfigure_CP_684_elements(27)); -- 
    cr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(27), ack => RPIPE_zeropad_input_pipe_336_inst_req_1); -- 
    -- CP-element group 28:  fork  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: 	32 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Sample/rr
      -- 
    ca_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_336_inst_ack_1, ack => testConfigure_CP_684_elements(28)); -- 
    rr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(28), ack => RPIPE_zeropad_input_pipe_342_inst_req_0); -- 
    -- CP-element group 29:  join  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (9) 
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/STORE_depth_high_338_Split/$entry
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/STORE_depth_high_338_Split/$exit
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/STORE_depth_high_338_Split/split_req
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/STORE_depth_high_338_Split/split_ack
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/word_access_start/$entry
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/word_access_start/word_0/$entry
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/word_access_start/word_0/rr
      -- 
    rr_1051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(29), ack => STORE_depth_high_338_store_0_req_0); -- 
    testConfigure_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(28) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (5) 
      -- CP-element group 30: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/word_access_start/$exit
      -- CP-element group 30: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/word_access_start/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/word_access_start/word_0/ra
      -- 
    ra_1052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_depth_high_338_store_0_ack_0, ack => testConfigure_CP_684_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	0 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	77 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/word_access_complete/$exit
      -- CP-element group 31: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/word_access_complete/word_0/$exit
      -- CP-element group 31: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/word_access_complete/word_0/ca
      -- 
    ca_1063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_depth_high_338_store_0_ack_1, ack => testConfigure_CP_684_elements(31)); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	28 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_update_start_
      -- CP-element group 32: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Update/cr
      -- 
    ra_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_342_inst_ack_0, ack => testConfigure_CP_684_elements(32)); -- 
    cr_1076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(32), ack => RPIPE_zeropad_input_pipe_342_inst_req_1); -- 
    -- CP-element group 33:  fork  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33: 	37 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Sample/rr
      -- 
    ca_1077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_342_inst_ack_1, ack => testConfigure_CP_684_elements(33)); -- 
    rr_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(33), ack => RPIPE_zeropad_input_pipe_348_inst_req_0); -- 
    -- CP-element group 34:  join  transition  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: 	0 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/STORE_pad_344_Split/$entry
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/STORE_pad_344_Split/$exit
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/STORE_pad_344_Split/split_req
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/STORE_pad_344_Split/split_ack
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/word_access_start/$entry
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/word_access_start/word_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/word_access_start/word_0/rr
      -- 
    rr_1098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(34), ack => STORE_pad_344_store_0_req_0); -- 
    testConfigure_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(33) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (5) 
      -- CP-element group 35: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/word_access_start/$exit
      -- CP-element group 35: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/word_access_start/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/word_access_start/word_0/ra
      -- 
    ra_1099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_pad_344_store_0_ack_0, ack => testConfigure_CP_684_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	77 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/word_access_complete/$exit
      -- CP-element group 36: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/word_access_complete/word_0/$exit
      -- CP-element group 36: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/word_access_complete/word_0/ca
      -- 
    ca_1110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_pad_344_store_0_ack_1, ack => testConfigure_CP_684_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	33 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_update_start_
      -- CP-element group 37: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Update/cr
      -- 
    ra_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_348_inst_ack_0, ack => testConfigure_CP_684_elements(37)); -- 
    cr_1123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(37), ack => RPIPE_zeropad_input_pipe_348_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	44 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Sample/rr
      -- 
    ca_1124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_348_inst_ack_1, ack => testConfigure_CP_684_elements(38)); -- 
    rr_1132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(38), ack => type_cast_352_inst_req_0); -- 
    rr_1196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(38), ack => RPIPE_zeropad_input_pipe_367_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Sample/ra
      -- 
    ra_1133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_352_inst_ack_0, ack => testConfigure_CP_684_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Update/ca
      -- 
    ca_1138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_352_inst_ack_1, ack => testConfigure_CP_684_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/ptr_deref_363_Split/$entry
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/ptr_deref_363_Split/$exit
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/ptr_deref_363_Split/split_req
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/ptr_deref_363_Split/split_ack
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/word_access_start/word_0/rr
      -- 
    rr_1176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(41), ack => ptr_deref_363_store_0_req_0); -- 
    testConfigure_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(40) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	75 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/word_access_start/$exit
      -- CP-element group 42: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/word_access_start/word_0/ra
      -- 
    ra_1177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_363_store_0_ack_0, ack => testConfigure_CP_684_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	0 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	77 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/word_access_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/word_access_complete/word_0/ca
      -- 
    ca_1188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_363_store_0_ack_1, ack => testConfigure_CP_684_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	38 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (6) 
      -- CP-element group 44: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_update_start_
      -- CP-element group 44: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Update/cr
      -- 
    ra_1197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_367_inst_ack_0, ack => testConfigure_CP_684_elements(44)); -- 
    cr_1201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(44), ack => RPIPE_zeropad_input_pipe_367_inst_req_1); -- 
    -- CP-element group 45:  fork  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: 	51 
    -- CP-element group 45:  members (9) 
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Sample/rr
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Sample/rr
      -- 
    ca_1202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_367_inst_ack_1, ack => testConfigure_CP_684_elements(45)); -- 
    rr_1274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(45), ack => RPIPE_zeropad_input_pipe_386_inst_req_0); -- 
    rr_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(45), ack => type_cast_371_inst_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Sample/ra
      -- 
    ra_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_0, ack => testConfigure_CP_684_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	0 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Update/ca
      -- 
    ca_1216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_1, ack => testConfigure_CP_684_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: 	75 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/ptr_deref_382_Split/$entry
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/ptr_deref_382_Split/$exit
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/ptr_deref_382_Split/split_req
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/ptr_deref_382_Split/split_ack
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/word_access_start/$entry
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/word_access_start/word_0/rr
      -- 
    rr_1254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(48), ack => ptr_deref_382_store_0_req_0); -- 
    testConfigure_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(47) & testConfigure_CP_684_elements(75) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	76 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/word_access_start/word_0/ra
      -- 
    ra_1255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_382_store_0_ack_0, ack => testConfigure_CP_684_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	0 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	77 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/word_access_complete/word_0/ca
      -- 
    ca_1266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_382_store_0_ack_1, ack => testConfigure_CP_684_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	45 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_update_start_
      -- CP-element group 51: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Update/cr
      -- 
    ra_1275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_386_inst_ack_0, ack => testConfigure_CP_684_elements(51)); -- 
    cr_1279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(51), ack => RPIPE_zeropad_input_pipe_386_inst_req_1); -- 
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Sample/rr
      -- 
    ca_1280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_386_inst_ack_1, ack => testConfigure_CP_684_elements(52)); -- 
    rr_1288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(52), ack => type_cast_390_inst_req_0); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Sample/ra
      -- 
    ra_1289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_390_inst_ack_0, ack => testConfigure_CP_684_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	0 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Update/ca
      -- 
    ca_1294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_390_inst_ack_1, ack => testConfigure_CP_684_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	76 
    -- CP-element group 55: 	54 
    -- CP-element group 55: 	0 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/ptr_deref_401_Split/$entry
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/ptr_deref_401_Split/$exit
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/ptr_deref_401_Split/split_req
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/ptr_deref_401_Split/split_ack
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/word_access_start/word_0/rr
      -- 
    rr_1332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(55), ack => ptr_deref_401_store_0_req_0); -- 
    testConfigure_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(76) & testConfigure_CP_684_elements(54) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/word_access_start/word_0/ra
      -- 
    ra_1333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_401_store_0_ack_0, ack => testConfigure_CP_684_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	77 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/word_access_complete/word_0/ca
      -- 
    ca_1344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_401_store_0_ack_1, ack => testConfigure_CP_684_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	72 
    -- CP-element group 58: 	0 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (5) 
      -- CP-element group 58: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/word_access_start/$entry
      -- CP-element group 58: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/word_access_start/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/word_access_start/word_0/rr
      -- 
    rr_1377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(58), ack => ptr_deref_414_load_0_req_0); -- 
    testConfigure_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(72) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/word_access_start/$exit
      -- CP-element group 59: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/word_access_start/word_0/$exit
      -- CP-element group 59: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/word_access_start/word_0/ra
      -- 
    ra_1378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_414_load_0_ack_0, ack => testConfigure_CP_684_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	67 
    -- CP-element group 60:  members (9) 
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/word_access_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/word_access_complete/word_0/$exit
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/word_access_complete/word_0/ca
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/ptr_deref_414_Merge/$entry
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/ptr_deref_414_Merge/$exit
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/ptr_deref_414_Merge/merge_req
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/ptr_deref_414_Merge/merge_ack
      -- 
    ca_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_414_load_0_ack_1, ack => testConfigure_CP_684_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	73 
    -- CP-element group 61: 	0 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/word_access_start/$entry
      -- CP-element group 61: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/word_access_start/word_0/rr
      -- 
    rr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(61), ack => ptr_deref_426_load_0_req_0); -- 
    testConfigure_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(73) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/word_access_start/$exit
      -- CP-element group 62: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/word_access_start/word_0/ra
      -- 
    ra_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_426_load_0_ack_0, ack => testConfigure_CP_684_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	0 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	67 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/word_access_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/word_access_complete/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/word_access_complete/word_0/ca
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/ptr_deref_426_Merge/$entry
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/ptr_deref_426_Merge/$exit
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/ptr_deref_426_Merge/merge_req
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/ptr_deref_426_Merge/merge_ack
      -- 
    ca_1439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_426_load_0_ack_1, ack => testConfigure_CP_684_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	74 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/word_access_start/$entry
      -- CP-element group 64: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/word_access_start/word_0/$entry
      -- CP-element group 64: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/word_access_start/word_0/rr
      -- 
    rr_1477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(64), ack => ptr_deref_438_load_0_req_0); -- 
    testConfigure_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(74) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/word_access_start/$exit
      -- CP-element group 65: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/word_access_start/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/word_access_start/word_0/ra
      -- 
    ra_1478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_438_load_0_ack_0, ack => testConfigure_CP_684_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	0 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (9) 
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/word_access_complete/$exit
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/word_access_complete/word_0/$exit
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/word_access_complete/word_0/ca
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/ptr_deref_438_Merge/$entry
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/ptr_deref_438_Merge/$exit
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/ptr_deref_438_Merge/merge_req
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/ptr_deref_438_Merge/merge_ack
      -- 
    ca_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_438_load_0_ack_1, ack => testConfigure_CP_684_elements(66)); -- 
    -- CP-element group 67:  join  transition  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	60 
    -- CP-element group 67: 	63 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Sample/rr
      -- 
    rr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(67), ack => type_cast_452_inst_req_0); -- 
    testConfigure_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(60) & testConfigure_CP_684_elements(63) & testConfigure_CP_684_elements(66);
      gj_testConfigure_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Sample/ra
      -- 
    ra_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_0, ack => testConfigure_CP_684_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	77 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Update/ca
      -- 
    ca_1508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_1, ack => testConfigure_CP_684_elements(69)); -- 
    -- CP-element group 70:  transition  delay-element  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	1 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	7 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_ptr_deref_303_delay
      -- 
    -- Element group testConfigure_CP_684_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(1), ack => testConfigure_CP_684_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  transition  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	8 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	14 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_ptr_deref_320_delay
      -- 
    -- Element group testConfigure_CP_684_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(8), ack => testConfigure_CP_684_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  delay-element  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	15 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	58 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_ptr_deref_414_delay
      -- 
    -- Element group testConfigure_CP_684_elements(72) is a control-delay.
    cp_element_72_delay: control_delay_element  generic map(name => " 72_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(15), ack => testConfigure_CP_684_elements(72), clk => clk, reset =>reset);
    -- CP-element group 73:  transition  delay-element  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	15 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	61 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_ptr_deref_426_delay
      -- 
    -- Element group testConfigure_CP_684_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(15), ack => testConfigure_CP_684_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  transition  delay-element  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	15 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	64 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_ptr_deref_438_delay
      -- 
    -- Element group testConfigure_CP_684_elements(74) is a control-delay.
    cp_element_74_delay: control_delay_element  generic map(name => " 74_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(15), ack => testConfigure_CP_684_elements(74), clk => clk, reset =>reset);
    -- CP-element group 75:  transition  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	42 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	48 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_ptr_deref_382_delay
      -- 
    -- Element group testConfigure_CP_684_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(42), ack => testConfigure_CP_684_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  transition  delay-element  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	49 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	55 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_ptr_deref_401_delay
      -- 
    -- Element group testConfigure_CP_684_elements(76) is a control-delay.
    cp_element_76_delay: control_delay_element  generic map(name => " 76_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(49), ack => testConfigure_CP_684_elements(76), clk => clk, reset =>reset);
    -- CP-element group 77:  branch  join  transition  place  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	9 
    -- CP-element group 77: 	21 
    -- CP-element group 77: 	57 
    -- CP-element group 77: 	26 
    -- CP-element group 77: 	69 
    -- CP-element group 77: 	31 
    -- CP-element group 77: 	36 
    -- CP-element group 77: 	50 
    -- CP-element group 77: 	16 
    -- CP-element group 77: 	43 
    -- CP-element group 77: 	2 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (10) 
      -- CP-element group 77: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465__exit__
      -- CP-element group 77: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/$exit
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466__entry__
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466_dead_link/$entry
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466_eval_test/$entry
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466_eval_test/$exit
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466_eval_test/branch_req
      -- CP-element group 77: 	 branch_block_stmt_277/R_cmp71_467_place
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466_if_link/$entry
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466_else_link/$entry
      -- 
    branch_req_1523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(77), ack => if_stmt_466_branch_req_0); -- 
    testConfigure_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(9) & testConfigure_CP_684_elements(21) & testConfigure_CP_684_elements(57) & testConfigure_CP_684_elements(26) & testConfigure_CP_684_elements(69) & testConfigure_CP_684_elements(31) & testConfigure_CP_684_elements(36) & testConfigure_CP_684_elements(50) & testConfigure_CP_684_elements(16) & testConfigure_CP_684_elements(43) & testConfigure_CP_684_elements(2);
      gj_testConfigure_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	132 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_277/if_stmt_466_if_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_277/if_stmt_466_if_link/if_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_277/entry_forx_xend
      -- CP-element group 78: 	 branch_block_stmt_277/entry_forx_xend_PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_277/entry_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_1528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_466_branch_ack_1, ack => testConfigure_CP_684_elements(78)); -- 
    -- CP-element group 79:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (18) 
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505__entry__
      -- CP-element group 79: 	 branch_block_stmt_277/merge_stmt_472__exit__
      -- CP-element group 79: 	 branch_block_stmt_277/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_277/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 79: 	 branch_block_stmt_277/merge_stmt_472_PhiReqMerge
      -- CP-element group 79: 	 branch_block_stmt_277/merge_stmt_472_PhiAck/$entry
      -- CP-element group 79: 	 branch_block_stmt_277/merge_stmt_472_PhiAck/$exit
      -- CP-element group 79: 	 branch_block_stmt_277/merge_stmt_472_PhiAck/dummy
      -- CP-element group 79: 	 branch_block_stmt_277/if_stmt_466_else_link/$exit
      -- CP-element group 79: 	 branch_block_stmt_277/if_stmt_466_else_link/else_choice_transition
      -- CP-element group 79: 	 branch_block_stmt_277/entry_bbx_xnph
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/$entry
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_update_start_
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Update/cr
      -- 
    else_choice_transition_1532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_466_branch_ack_0, ack => testConfigure_CP_684_elements(79)); -- 
    rr_1545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(79), ack => type_cast_485_inst_req_0); -- 
    cr_1550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(79), ack => type_cast_485_inst_req_1); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Sample/ra
      -- 
    ra_1546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_485_inst_ack_0, ack => testConfigure_CP_684_elements(80)); -- 
    -- CP-element group 81:  transition  place  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	126 
    -- CP-element group 81:  members (9) 
      -- CP-element group 81: 	 branch_block_stmt_277/bbx_xnph_forx_xbody
      -- CP-element group 81: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505__exit__
      -- CP-element group 81: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 81: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/$entry
      -- CP-element group 81: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/phi_stmt_508/$entry
      -- CP-element group 81: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/$exit
      -- CP-element group 81: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Update/ca
      -- 
    ca_1551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_485_inst_ack_1, ack => testConfigure_CP_684_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	131 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	121 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_sample_complete
      -- CP-element group 82: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Sample/ack
      -- 
    ack_1580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_520_index_offset_ack_0, ack => testConfigure_CP_684_elements(82)); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	131 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (11) 
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_request/$entry
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_base_plus_offset/$entry
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_request/req
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Update/ack
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_base_plus_offset/$exit
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_base_plus_offset/sum_rename_req
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_base_plus_offset/sum_rename_ack
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_root_address_calculated
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_offset_calculated
      -- 
    ack_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_520_index_offset_ack_1, ack => testConfigure_CP_684_elements(83)); -- 
    req_1594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(83), ack => addr_of_521_final_reg_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_request/$exit
      -- CP-element group 84: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_request/ack
      -- CP-element group 84: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_sample_completed_
      -- 
    ack_1595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_521_final_reg_ack_0, ack => testConfigure_CP_684_elements(84)); -- 
    -- CP-element group 85:  fork  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	131 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (19) 
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_word_addrgen/$entry
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_addr_resize/$exit
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_word_addrgen/$exit
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_addr_resize/$entry
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_address_resized
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_plus_offset/sum_rename_ack
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_complete/$exit
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_complete/ack
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_word_addrgen/root_register_req
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_word_addrgen/root_register_ack
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_addr_resize/base_resize_req
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_addr_resize/base_resize_ack
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_plus_offset/sum_rename_req
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_plus_offset/$exit
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_plus_offset/$entry
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_root_address_calculated
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_word_address_calculated
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_address_calculated
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_update_completed_
      -- 
    ack_1600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_521_final_reg_ack_1, ack => testConfigure_CP_684_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	131 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Update/cr
      -- CP-element group 86: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_update_start_
      -- 
    ra_1609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_524_inst_ack_0, ack => testConfigure_CP_684_elements(86)); -- 
    cr_1613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(86), ack => RPIPE_zeropad_input_pipe_524_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_update_completed_
      -- 
    ca_1614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_524_inst_ack_1, ack => testConfigure_CP_684_elements(87)); -- 
    rr_1622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(87), ack => type_cast_528_inst_req_0); -- 
    rr_1636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(87), ack => RPIPE_zeropad_input_pipe_537_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Sample/ra
      -- CP-element group 88: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_sample_completed_
      -- 
    ra_1623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_528_inst_ack_0, ack => testConfigure_CP_684_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	131 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Update/ca
      -- CP-element group 89: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_update_completed_
      -- 
    ca_1628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_528_inst_ack_1, ack => testConfigure_CP_684_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_update_start_
      -- CP-element group 90: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Update/cr
      -- 
    ra_1637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_537_inst_ack_0, ack => testConfigure_CP_684_elements(90)); -- 
    cr_1641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(90), ack => RPIPE_zeropad_input_pipe_537_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Sample/$entry
      -- 
    ca_1642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_537_inst_ack_1, ack => testConfigure_CP_684_elements(91)); -- 
    rr_1650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(91), ack => type_cast_541_inst_req_0); -- 
    rr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(91), ack => RPIPE_zeropad_input_pipe_555_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Sample/ra
      -- 
    ra_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_541_inst_ack_0, ack => testConfigure_CP_684_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	131 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Update/ca
      -- 
    ca_1656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_541_inst_ack_1, ack => testConfigure_CP_684_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_update_start_
      -- 
    ra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_555_inst_ack_0, ack => testConfigure_CP_684_elements(94)); -- 
    cr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(94), ack => RPIPE_zeropad_input_pipe_555_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_sample_start_
      -- 
    ca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_555_inst_ack_1, ack => testConfigure_CP_684_elements(95)); -- 
    rr_1678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(95), ack => type_cast_559_inst_req_0); -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(95), ack => RPIPE_zeropad_input_pipe_573_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Sample/ra
      -- 
    ra_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_559_inst_ack_0, ack => testConfigure_CP_684_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	131 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Update/$exit
      -- 
    ca_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_559_inst_ack_1, ack => testConfigure_CP_684_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_update_start_
      -- CP-element group 98: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_sample_completed_
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_573_inst_ack_0, ack => testConfigure_CP_684_elements(98)); -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(98), ack => RPIPE_zeropad_input_pipe_573_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_update_completed_
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_573_inst_ack_1, ack => testConfigure_CP_684_elements(99)); -- 
    rr_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(99), ack => type_cast_577_inst_req_0); -- 
    rr_1720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(99), ack => RPIPE_zeropad_input_pipe_591_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_sample_completed_
      -- 
    ra_1707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_0, ack => testConfigure_CP_684_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	131 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Update/ca
      -- CP-element group 101: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_update_completed_
      -- 
    ca_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_1, ack => testConfigure_CP_684_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_update_start_
      -- CP-element group 102: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_sample_completed_
      -- 
    ra_1721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_591_inst_ack_0, ack => testConfigure_CP_684_elements(102)); -- 
    cr_1725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(102), ack => RPIPE_zeropad_input_pipe_591_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_update_completed_
      -- 
    ca_1726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_591_inst_ack_1, ack => testConfigure_CP_684_elements(103)); -- 
    rr_1734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(103), ack => type_cast_595_inst_req_0); -- 
    rr_1748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(103), ack => RPIPE_zeropad_input_pipe_609_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_sample_completed_
      -- 
    ra_1735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_595_inst_ack_0, ack => testConfigure_CP_684_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	131 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_update_completed_
      -- 
    ca_1740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_595_inst_ack_1, ack => testConfigure_CP_684_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Update/cr
      -- CP-element group 106: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_update_start_
      -- CP-element group 106: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Update/$entry
      -- 
    ra_1749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_609_inst_ack_0, ack => testConfigure_CP_684_elements(106)); -- 
    cr_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(106), ack => RPIPE_zeropad_input_pipe_609_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Sample/rr
      -- 
    ca_1754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_609_inst_ack_1, ack => testConfigure_CP_684_elements(107)); -- 
    rr_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(107), ack => type_cast_613_inst_req_0); -- 
    rr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(107), ack => RPIPE_zeropad_input_pipe_627_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Sample/ra
      -- 
    ra_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_613_inst_ack_0, ack => testConfigure_CP_684_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	131 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Update/ca
      -- 
    ca_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_613_inst_ack_1, ack => testConfigure_CP_684_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_update_start_
      -- CP-element group 110: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Update/cr
      -- 
    ra_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_627_inst_ack_0, ack => testConfigure_CP_684_elements(110)); -- 
    cr_1781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(110), ack => RPIPE_zeropad_input_pipe_627_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Sample/$entry
      -- 
    ca_1782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_627_inst_ack_1, ack => testConfigure_CP_684_elements(111)); -- 
    rr_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(111), ack => type_cast_631_inst_req_0); -- 
    rr_1804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(111), ack => RPIPE_zeropad_input_pipe_645_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Sample/ra
      -- CP-element group 112: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_sample_completed_
      -- 
    ra_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_631_inst_ack_0, ack => testConfigure_CP_684_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	131 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Update/ca
      -- CP-element group 113: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_update_completed_
      -- 
    ca_1796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_631_inst_ack_1, ack => testConfigure_CP_684_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_update_start_
      -- CP-element group 114: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Sample/$exit
      -- 
    ra_1805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_645_inst_ack_0, ack => testConfigure_CP_684_elements(114)); -- 
    cr_1809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(114), ack => RPIPE_zeropad_input_pipe_645_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Update/$exit
      -- 
    ca_1810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_645_inst_ack_1, ack => testConfigure_CP_684_elements(115)); -- 
    rr_1818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(115), ack => type_cast_649_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_sample_completed_
      -- 
    ra_1819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_0, ack => testConfigure_CP_684_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	131 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_update_completed_
      -- 
    ca_1824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_1, ack => testConfigure_CP_684_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (9) 
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/ptr_deref_657_Split/split_req
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/ptr_deref_657_Split/split_ack
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/word_access_start/$entry
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/word_access_start/word_0/$entry
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/ptr_deref_657_Split/$exit
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/ptr_deref_657_Split/$entry
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/word_access_start/word_0/rr
      -- 
    rr_1862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(118), ack => ptr_deref_657_store_0_req_0); -- 
    testConfigure_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(85) & testConfigure_CP_684_elements(89) & testConfigure_CP_684_elements(93) & testConfigure_CP_684_elements(97) & testConfigure_CP_684_elements(101) & testConfigure_CP_684_elements(105) & testConfigure_CP_684_elements(109) & testConfigure_CP_684_elements(113) & testConfigure_CP_684_elements(117);
      gj_testConfigure_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/word_access_start/$exit
      -- CP-element group 119: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/word_access_start/word_0/$exit
      -- CP-element group 119: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/word_access_start/word_0/ra
      -- 
    ra_1863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_657_store_0_ack_0, ack => testConfigure_CP_684_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	131 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/word_access_complete/word_0/ca
      -- CP-element group 120: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/word_access_complete/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/word_access_complete/$exit
      -- CP-element group 120: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/$exit
      -- 
    ca_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_657_store_0_ack_1, ack => testConfigure_CP_684_elements(120)); -- 
    -- CP-element group 121:  branch  join  transition  place  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	82 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (10) 
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671__entry__
      -- CP-element group 121: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670__exit__
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671_if_link/$entry
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671_else_link/$entry
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671_eval_test/branch_req
      -- CP-element group 121: 	 branch_block_stmt_277/R_exitcond7_672_place
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671_dead_link/$entry
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671_eval_test/$entry
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671_eval_test/$exit
      -- CP-element group 121: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/$exit
      -- 
    branch_req_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(121), ack => if_stmt_671_branch_req_0); -- 
    testConfigure_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(82) & testConfigure_CP_684_elements(120);
      gj_testConfigure_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  merge  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	132 
    -- CP-element group 122:  members (13) 
      -- CP-element group 122: 	 branch_block_stmt_277/forx_xendx_xloopexit_forx_xend
      -- CP-element group 122: 	 branch_block_stmt_277/merge_stmt_677__exit__
      -- CP-element group 122: 	 branch_block_stmt_277/if_stmt_671_if_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_277/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 122: 	 branch_block_stmt_277/if_stmt_671_if_link/if_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_277/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_277/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 122: 	 branch_block_stmt_277/merge_stmt_677_PhiReqMerge
      -- CP-element group 122: 	 branch_block_stmt_277/merge_stmt_677_PhiAck/$entry
      -- CP-element group 122: 	 branch_block_stmt_277/merge_stmt_677_PhiAck/$exit
      -- CP-element group 122: 	 branch_block_stmt_277/merge_stmt_677_PhiAck/dummy
      -- CP-element group 122: 	 branch_block_stmt_277/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_277/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_1887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_671_branch_ack_1, ack => testConfigure_CP_684_elements(122)); -- 
    -- CP-element group 123:  fork  transition  place  input  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	127 
    -- CP-element group 123: 	128 
    -- CP-element group 123:  members (12) 
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody
      -- CP-element group 123: 	 branch_block_stmt_277/if_stmt_671_else_link/$exit
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Update/cr
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Sample/rr
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/if_stmt_671_else_link/else_choice_transition
      -- 
    else_choice_transition_1891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_671_branch_ack_0, ack => testConfigure_CP_684_elements(123)); -- 
    cr_1957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(123), ack => type_cast_514_inst_req_1); -- 
    rr_1952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(123), ack => type_cast_514_inst_req_0); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	132 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Sample/ra
      -- 
    ra_1905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_682_inst_ack_0, ack => testConfigure_CP_684_elements(124)); -- 
    -- CP-element group 125:  transition  place  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	132 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (16) 
      -- CP-element group 125: 	 branch_block_stmt_277/branch_block_stmt_277__exit__
      -- CP-element group 125: 	 branch_block_stmt_277/merge_stmt_685__exit__
      -- CP-element group 125: 	 branch_block_stmt_277/return__
      -- CP-element group 125: 	 branch_block_stmt_277/assign_stmt_683__exit__
      -- CP-element group 125: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_277/$exit
      -- CP-element group 125: 	 $exit
      -- CP-element group 125: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_277/assign_stmt_683/$exit
      -- CP-element group 125: 	 branch_block_stmt_277/return___PhiReq/$entry
      -- CP-element group 125: 	 branch_block_stmt_277/return___PhiReq/$exit
      -- CP-element group 125: 	 branch_block_stmt_277/merge_stmt_685_PhiReqMerge
      -- CP-element group 125: 	 branch_block_stmt_277/merge_stmt_685_PhiAck/$entry
      -- CP-element group 125: 	 branch_block_stmt_277/merge_stmt_685_PhiAck/$exit
      -- CP-element group 125: 	 branch_block_stmt_277/merge_stmt_685_PhiAck/dummy
      -- 
    ca_1910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_682_inst_ack_1, ack => testConfigure_CP_684_elements(125)); -- 
    -- CP-element group 126:  transition  output  delay-element  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	81 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	130 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_req
      -- CP-element group 126: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 126: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/$exit
      -- CP-element group 126: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_512_konst_delay_trans
      -- CP-element group 126: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/phi_stmt_508/$exit
      -- 
    phi_stmt_508_req_1933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_508_req_1933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(126), ack => phi_stmt_508_req_0); -- 
    -- Element group testConfigure_CP_684_elements(126) is a control-delay.
    cp_element_126_delay: control_delay_element  generic map(name => " 126_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(81), ack => testConfigure_CP_684_elements(126), clk => clk, reset =>reset);
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	123 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Sample/ra
      -- 
    ra_1953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_514_inst_ack_0, ack => testConfigure_CP_684_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	123 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Update/ca
      -- CP-element group 128: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Update/$exit
      -- 
    ca_1958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_514_inst_ack_1, ack => testConfigure_CP_684_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 129: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/$exit
      -- CP-element group 129: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/$exit
      -- CP-element group 129: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_req
      -- CP-element group 129: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/$exit
      -- CP-element group 129: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/$exit
      -- 
    phi_stmt_508_req_1959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_508_req_1959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(129), ack => phi_stmt_508_req_1); -- 
    testConfigure_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(127) & testConfigure_CP_684_elements(128);
      gj_testConfigure_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  merge  transition  place  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	126 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_277/merge_stmt_507_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_277/merge_stmt_507_PhiAck/$entry
      -- 
    testConfigure_CP_684_elements(130) <= OrReduce(testConfigure_CP_684_elements(126) & testConfigure_CP_684_elements(129));
    -- CP-element group 131:  fork  transition  place  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	82 
    -- CP-element group 131: 	83 
    -- CP-element group 131: 	85 
    -- CP-element group 131: 	86 
    -- CP-element group 131: 	89 
    -- CP-element group 131: 	93 
    -- CP-element group 131: 	97 
    -- CP-element group 131: 	101 
    -- CP-element group 131: 	105 
    -- CP-element group 131: 	109 
    -- CP-element group 131: 	113 
    -- CP-element group 131: 	117 
    -- CP-element group 131: 	120 
    -- CP-element group 131:  members (56) 
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_resize_1/index_resize_ack
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_update_start
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_scale_1/$exit
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670__entry__
      -- CP-element group 131: 	 branch_block_stmt_277/merge_stmt_507__exit__
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_scale_1/scale_rename_req
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Sample/req
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_scale_1/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_scale_1/scale_rename_ack
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_complete/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_complete/req
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Update/req
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/word_access_complete/word_0/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/word_access_complete/word_0/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/word_access_complete/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_resize_1/index_resize_req
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_resize_1/$exit
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_resize_1/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_computed_1
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_resized_1
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_scaled_1
      -- CP-element group 131: 	 branch_block_stmt_277/merge_stmt_507_PhiAck/$exit
      -- CP-element group 131: 	 branch_block_stmt_277/merge_stmt_507_PhiAck/phi_stmt_508_ack
      -- 
    phi_stmt_508_ack_1964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_508_ack_0, ack => testConfigure_CP_684_elements(131)); -- 
    cr_1739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_595_inst_req_1); -- 
    cr_1627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_528_inst_req_1); -- 
    req_1579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => array_obj_ref_520_index_offset_req_0); -- 
    cr_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_613_inst_req_1); -- 
    cr_1795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_631_inst_req_1); -- 
    req_1599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => addr_of_521_final_reg_req_1); -- 
    req_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => array_obj_ref_520_index_offset_req_1); -- 
    cr_1655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_541_inst_req_1); -- 
    cr_1823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_649_inst_req_1); -- 
    cr_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => ptr_deref_657_store_0_req_1); -- 
    cr_1711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_577_inst_req_1); -- 
    rr_1608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => RPIPE_zeropad_input_pipe_524_inst_req_0); -- 
    cr_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_559_inst_req_1); -- 
    -- CP-element group 132:  merge  fork  transition  place  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	78 
    -- CP-element group 132: 	122 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	124 
    -- CP-element group 132: 	125 
    -- CP-element group 132:  members (13) 
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683__entry__
      -- CP-element group 132: 	 branch_block_stmt_277/merge_stmt_679__exit__
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_update_start_
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/$entry
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_277/merge_stmt_679_PhiReqMerge
      -- CP-element group 132: 	 branch_block_stmt_277/merge_stmt_679_PhiAck/$entry
      -- CP-element group 132: 	 branch_block_stmt_277/merge_stmt_679_PhiAck/$exit
      -- CP-element group 132: 	 branch_block_stmt_277/merge_stmt_679_PhiAck/dummy
      -- 
    rr_1904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(132), ack => type_cast_682_inst_req_0); -- 
    cr_1909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(132), ack => type_cast_682_inst_req_1); -- 
    testConfigure_CP_684_elements(132) <= OrReduce(testConfigure_CP_684_elements(78) & testConfigure_CP_684_elements(122));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_519_resized : std_logic_vector(13 downto 0);
    signal R_indvar_519_scaled : std_logic_vector(13 downto 0);
    signal STORE_col_high_332_data_0 : std_logic_vector(7 downto 0);
    signal STORE_col_high_332_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_depth_high_338_data_0 : std_logic_vector(7 downto 0);
    signal STORE_depth_high_338_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_pad_344_data_0 : std_logic_vector(7 downto 0);
    signal STORE_pad_344_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_row_high_326_data_0 : std_logic_vector(7 downto 0);
    signal STORE_row_high_326_word_address_0 : std_logic_vector(0 downto 0);
    signal add33_565 : std_logic_vector(63 downto 0);
    signal add39_583 : std_logic_vector(63 downto 0);
    signal add45_601 : std_logic_vector(63 downto 0);
    signal add51_619 : std_logic_vector(63 downto 0);
    signal add57_637 : std_logic_vector(63 downto 0);
    signal add63_655 : std_logic_vector(63 downto 0);
    signal add_547 : std_logic_vector(63 downto 0);
    signal array_obj_ref_520_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_520_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_520_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_520_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_520_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_520_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_522 : std_logic_vector(31 downto 0);
    signal call11_387 : std_logic_vector(7 downto 0);
    signal call1_308 : std_logic_vector(7 downto 0);
    signal call22_525 : std_logic_vector(7 downto 0);
    signal call25_538 : std_logic_vector(7 downto 0);
    signal call30_556 : std_logic_vector(7 downto 0);
    signal call36_574 : std_logic_vector(7 downto 0);
    signal call3_325 : std_logic_vector(7 downto 0);
    signal call42_592 : std_logic_vector(7 downto 0);
    signal call48_610 : std_logic_vector(7 downto 0);
    signal call4_331 : std_logic_vector(7 downto 0);
    signal call54_628 : std_logic_vector(7 downto 0);
    signal call5_337 : std_logic_vector(7 downto 0);
    signal call60_646 : std_logic_vector(7 downto 0);
    signal call6_343 : std_logic_vector(7 downto 0);
    signal call7_349 : std_logic_vector(7 downto 0);
    signal call9_368 : std_logic_vector(7 downto 0);
    signal call_291 : std_logic_vector(7 downto 0);
    signal cmp71_465 : std_logic_vector(0 downto 0);
    signal conv10_372 : std_logic_vector(31 downto 0);
    signal conv12_391 : std_logic_vector(31 downto 0);
    signal conv16_453 : std_logic_vector(63 downto 0);
    signal conv23_529 : std_logic_vector(63 downto 0);
    signal conv27_542 : std_logic_vector(63 downto 0);
    signal conv2_312 : std_logic_vector(31 downto 0);
    signal conv32_560 : std_logic_vector(63 downto 0);
    signal conv38_578 : std_logic_vector(63 downto 0);
    signal conv44_596 : std_logic_vector(63 downto 0);
    signal conv50_614 : std_logic_vector(63 downto 0);
    signal conv56_632 : std_logic_vector(63 downto 0);
    signal conv62_650 : std_logic_vector(63 downto 0);
    signal conv8_353 : std_logic_vector(31 downto 0);
    signal conv_295 : std_logic_vector(31 downto 0);
    signal exitcond7_670 : std_logic_vector(0 downto 0);
    signal iNsTr_0_283 : std_logic_vector(31 downto 0);
    signal iNsTr_17_361 : std_logic_vector(31 downto 0);
    signal iNsTr_20_380 : std_logic_vector(31 downto 0);
    signal iNsTr_23_399 : std_logic_vector(31 downto 0);
    signal iNsTr_25_411 : std_logic_vector(31 downto 0);
    signal iNsTr_26_423 : std_logic_vector(31 downto 0);
    signal iNsTr_27_435 : std_logic_vector(31 downto 0);
    signal iNsTr_3_301 : std_logic_vector(31 downto 0);
    signal iNsTr_6_318 : std_logic_vector(31 downto 0);
    signal indvar_508 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_665 : std_logic_vector(63 downto 0);
    signal mul15_449 : std_logic_vector(31 downto 0);
    signal mul_444 : std_logic_vector(31 downto 0);
    signal ptr_deref_285_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_285_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_285_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_285_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_285_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_285_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_303_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_303_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_303_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_303_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_303_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_303_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_320_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_320_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_320_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_320_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_320_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_320_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_363_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_363_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_363_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_363_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_363_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_363_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_382_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_382_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_382_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_382_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_382_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_382_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_401_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_401_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_401_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_401_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_401_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_401_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_414_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_414_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_414_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_414_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_414_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_426_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_426_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_426_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_426_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_426_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_438_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_438_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_438_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_438_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_438_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_657_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_657_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_657_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_657_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_657_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_657_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl29_553 : std_logic_vector(63 downto 0);
    signal shl35_571 : std_logic_vector(63 downto 0);
    signal shl41_589 : std_logic_vector(63 downto 0);
    signal shl47_607 : std_logic_vector(63 downto 0);
    signal shl53_625 : std_logic_vector(63 downto 0);
    signal shl59_643 : std_logic_vector(63 downto 0);
    signal shl_535 : std_logic_vector(63 downto 0);
    signal shr70x_xmask_459 : std_logic_vector(63 downto 0);
    signal tmp13_427 : std_logic_vector(31 downto 0);
    signal tmp14_439 : std_logic_vector(31 downto 0);
    signal tmp1_477 : std_logic_vector(31 downto 0);
    signal tmp2_482 : std_logic_vector(31 downto 0);
    signal tmp3_486 : std_logic_vector(63 downto 0);
    signal tmp4_492 : std_logic_vector(63 downto 0);
    signal tmp5_498 : std_logic_vector(0 downto 0);
    signal tmp_415 : std_logic_vector(31 downto 0);
    signal type_cast_287_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_457_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_463_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_490_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_496_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_503_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_512_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_514_wire : std_logic_vector(63 downto 0);
    signal type_cast_533_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_551_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_569_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_587_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_605_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_623_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_641_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_663_wire_constant : std_logic_vector(63 downto 0);
    signal umax6_505 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_col_high_332_word_address_0 <= "0";
    STORE_depth_high_338_word_address_0 <= "0";
    STORE_pad_344_word_address_0 <= "0";
    STORE_row_high_326_word_address_0 <= "0";
    array_obj_ref_520_constant_part_of_offset <= "00000000000000";
    array_obj_ref_520_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_520_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_520_resized_base_address <= "00000000000000";
    iNsTr_0_283 <= "00000000000000000000000000000000";
    iNsTr_17_361 <= "00000000000000000000000000000011";
    iNsTr_20_380 <= "00000000000000000000000000000100";
    iNsTr_23_399 <= "00000000000000000000000000000101";
    iNsTr_25_411 <= "00000000000000000000000000000011";
    iNsTr_26_423 <= "00000000000000000000000000000100";
    iNsTr_27_435 <= "00000000000000000000000000000101";
    iNsTr_3_301 <= "00000000000000000000000000000001";
    iNsTr_6_318 <= "00000000000000000000000000000010";
    ptr_deref_285_word_offset_0 <= "0000000";
    ptr_deref_303_word_offset_0 <= "0000000";
    ptr_deref_320_word_offset_0 <= "0000000";
    ptr_deref_363_word_offset_0 <= "0000000";
    ptr_deref_382_word_offset_0 <= "0000000";
    ptr_deref_401_word_offset_0 <= "0000000";
    ptr_deref_414_word_offset_0 <= "0000000";
    ptr_deref_426_word_offset_0 <= "0000000";
    ptr_deref_438_word_offset_0 <= "0000000";
    ptr_deref_657_word_offset_0 <= "00000000000000";
    type_cast_287_wire_constant <= "00000000000000000000000000000101";
    type_cast_457_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_463_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_490_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_496_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_503_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_512_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_533_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_551_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_569_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_587_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_605_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_623_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_641_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_663_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_508: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_512_wire_constant & type_cast_514_wire;
      req <= phi_stmt_508_req_0 & phi_stmt_508_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_508",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_508_ack_0,
          idata => idata,
          odata => indvar_508,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_508
    -- flow-through select operator MUX_504_inst
    umax6_505 <= tmp4_492 when (tmp5_498(0) /=  '0') else type_cast_503_wire_constant;
    addr_of_521_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_521_final_reg_req_0;
      addr_of_521_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_521_final_reg_req_1;
      addr_of_521_final_reg_ack_1<= rack(0);
      addr_of_521_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_521_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_520_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_522,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_294_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_294_inst_req_0;
      type_cast_294_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_294_inst_req_1;
      type_cast_294_inst_ack_1<= rack(0);
      type_cast_294_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_294_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_291,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_295,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_311_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_311_inst_req_0;
      type_cast_311_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_311_inst_req_1;
      type_cast_311_inst_ack_1<= rack(0);
      type_cast_311_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_311_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_308,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_312,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_352_inst_req_0;
      type_cast_352_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_352_inst_req_1;
      type_cast_352_inst_ack_1<= rack(0);
      type_cast_352_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_352_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call7_349,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_353,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_371_inst_req_0;
      type_cast_371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_371_inst_req_1;
      type_cast_371_inst_ack_1<= rack(0);
      type_cast_371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call9_368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10_372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_390_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_390_inst_req_0;
      type_cast_390_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_390_inst_req_1;
      type_cast_390_inst_ack_1<= rack(0);
      type_cast_390_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_390_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_387,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_391,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_452_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_452_inst_req_0;
      type_cast_452_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_452_inst_req_1;
      type_cast_452_inst_ack_1<= rack(0);
      type_cast_452_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_452_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul15_449,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_453,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_485_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_485_inst_req_0;
      type_cast_485_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_485_inst_req_1;
      type_cast_485_inst_ack_1<= rack(0);
      type_cast_485_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_485_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp2_482,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_486,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_514_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_514_inst_req_0;
      type_cast_514_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_514_inst_req_1;
      type_cast_514_inst_ack_1<= rack(0);
      type_cast_514_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_514_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_665,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_514_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_528_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_528_inst_req_0;
      type_cast_528_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_528_inst_req_1;
      type_cast_528_inst_ack_1<= rack(0);
      type_cast_528_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_528_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_525,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_529,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_541_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_541_inst_req_0;
      type_cast_541_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_541_inst_req_1;
      type_cast_541_inst_ack_1<= rack(0);
      type_cast_541_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_541_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call25_538,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_542,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_559_inst_req_0;
      type_cast_559_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_559_inst_req_1;
      type_cast_559_inst_ack_1<= rack(0);
      type_cast_559_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_559_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call30_556,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_560,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_577_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_577_inst_req_0;
      type_cast_577_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_577_inst_req_1;
      type_cast_577_inst_ack_1<= rack(0);
      type_cast_577_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_577_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_574,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_578,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_595_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_595_inst_req_0;
      type_cast_595_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_595_inst_req_1;
      type_cast_595_inst_ack_1<= rack(0);
      type_cast_595_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_595_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call42_592,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_596,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_613_inst_req_0;
      type_cast_613_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_613_inst_req_1;
      type_cast_613_inst_ack_1<= rack(0);
      type_cast_613_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_613_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call48_610,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_614,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_631_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_631_inst_req_0;
      type_cast_631_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_631_inst_req_1;
      type_cast_631_inst_ack_1<= rack(0);
      type_cast_631_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_631_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call54_628,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_632,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_649_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_649_inst_req_0;
      type_cast_649_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_649_inst_req_1;
      type_cast_649_inst_ack_1<= rack(0);
      type_cast_649_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_649_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call60_646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_650,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_682_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_682_inst_req_0;
      type_cast_682_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_682_inst_req_1;
      type_cast_682_inst_ack_1<= rack(0);
      type_cast_682_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_682_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul15_449,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ret_val_x_x_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_col_high_332_gather_scatter
    process(call4_331) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call4_331;
      ov(7 downto 0) := iv;
      STORE_col_high_332_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_depth_high_338_gather_scatter
    process(call5_337) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call5_337;
      ov(7 downto 0) := iv;
      STORE_depth_high_338_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_pad_344_gather_scatter
    process(call6_343) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call6_343;
      ov(7 downto 0) := iv;
      STORE_pad_344_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_row_high_326_gather_scatter
    process(call3_325) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call3_325;
      ov(7 downto 0) := iv;
      STORE_row_high_326_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_520_index_1_rename
    process(R_indvar_519_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_519_resized;
      ov(13 downto 0) := iv;
      R_indvar_519_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_520_index_1_resize
    process(indvar_508) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_508;
      ov := iv(13 downto 0);
      R_indvar_519_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_520_root_address_inst
    process(array_obj_ref_520_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_520_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_520_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_285_addr_0
    process(ptr_deref_285_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_285_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_285_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_285_base_resize
    process(iNsTr_0_283) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_283;
      ov := iv(6 downto 0);
      ptr_deref_285_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_285_gather_scatter
    process(type_cast_287_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_287_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_285_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_285_root_address_inst
    process(ptr_deref_285_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_285_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_285_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_303_addr_0
    process(ptr_deref_303_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_303_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_303_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_303_base_resize
    process(iNsTr_3_301) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_301;
      ov := iv(6 downto 0);
      ptr_deref_303_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_303_gather_scatter
    process(conv_295) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_295;
      ov(31 downto 0) := iv;
      ptr_deref_303_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_303_root_address_inst
    process(ptr_deref_303_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_303_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_303_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_320_addr_0
    process(ptr_deref_320_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_320_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_320_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_320_base_resize
    process(iNsTr_6_318) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_318;
      ov := iv(6 downto 0);
      ptr_deref_320_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_320_gather_scatter
    process(conv2_312) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv2_312;
      ov(31 downto 0) := iv;
      ptr_deref_320_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_320_root_address_inst
    process(ptr_deref_320_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_320_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_320_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_363_addr_0
    process(ptr_deref_363_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_363_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_363_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_363_base_resize
    process(iNsTr_17_361) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_17_361;
      ov := iv(6 downto 0);
      ptr_deref_363_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_363_gather_scatter
    process(conv8_353) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv8_353;
      ov(31 downto 0) := iv;
      ptr_deref_363_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_363_root_address_inst
    process(ptr_deref_363_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_363_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_363_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_382_addr_0
    process(ptr_deref_382_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_382_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_382_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_382_base_resize
    process(iNsTr_20_380) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_20_380;
      ov := iv(6 downto 0);
      ptr_deref_382_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_382_gather_scatter
    process(conv10_372) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv10_372;
      ov(31 downto 0) := iv;
      ptr_deref_382_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_382_root_address_inst
    process(ptr_deref_382_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_382_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_382_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_401_addr_0
    process(ptr_deref_401_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_401_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_401_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_401_base_resize
    process(iNsTr_23_399) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_23_399;
      ov := iv(6 downto 0);
      ptr_deref_401_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_401_gather_scatter
    process(conv12_391) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv12_391;
      ov(31 downto 0) := iv;
      ptr_deref_401_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_401_root_address_inst
    process(ptr_deref_401_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_401_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_401_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_414_addr_0
    process(ptr_deref_414_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_414_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_414_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_414_base_resize
    process(iNsTr_25_411) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_25_411;
      ov := iv(6 downto 0);
      ptr_deref_414_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_414_gather_scatter
    process(ptr_deref_414_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_414_data_0;
      ov(31 downto 0) := iv;
      tmp_415 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_414_root_address_inst
    process(ptr_deref_414_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_414_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_414_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_addr_0
    process(ptr_deref_426_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_426_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_426_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_base_resize
    process(iNsTr_26_423) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_26_423;
      ov := iv(6 downto 0);
      ptr_deref_426_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_gather_scatter
    process(ptr_deref_426_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_426_data_0;
      ov(31 downto 0) := iv;
      tmp13_427 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_root_address_inst
    process(ptr_deref_426_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_426_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_426_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_438_addr_0
    process(ptr_deref_438_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_438_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_438_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_438_base_resize
    process(iNsTr_27_435) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_27_435;
      ov := iv(6 downto 0);
      ptr_deref_438_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_438_gather_scatter
    process(ptr_deref_438_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_438_data_0;
      ov(31 downto 0) := iv;
      tmp14_439 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_438_root_address_inst
    process(ptr_deref_438_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_438_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_438_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_657_addr_0
    process(ptr_deref_657_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_657_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_657_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_657_base_resize
    process(arrayidx_522) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_522;
      ov := iv(13 downto 0);
      ptr_deref_657_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_657_gather_scatter
    process(add63_655) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add63_655;
      ov(63 downto 0) := iv;
      ptr_deref_657_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_657_root_address_inst
    process(ptr_deref_657_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_657_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_657_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_466_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp71_465;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_466_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_466_branch_req_0,
          ack0 => if_stmt_466_branch_ack_0,
          ack1 => if_stmt_466_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_671_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond7_670;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_671_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_671_branch_req_0,
          ack0 => if_stmt_671_branch_ack_0,
          ack1 => if_stmt_671_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_664_inst
    process(indvar_508) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_508, type_cast_663_wire_constant, tmp_var);
      indvarx_xnext_665 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_458_inst
    process(conv16_453) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv16_453, type_cast_457_wire_constant, tmp_var);
      shr70x_xmask_459 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_464_inst
    process(shr70x_xmask_459) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr70x_xmask_459, type_cast_463_wire_constant, tmp_var);
      cmp71_465 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_669_inst
    process(indvarx_xnext_665, umax6_505) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_665, umax6_505, tmp_var);
      exitcond7_670 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_491_inst
    process(tmp3_486) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp3_486, type_cast_490_wire_constant, tmp_var);
      tmp4_492 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_443_inst
    process(tmp13_427, tmp_415) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp13_427, tmp_415, tmp_var);
      mul_444 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_448_inst
    process(mul_444, tmp14_439) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_444, tmp14_439, tmp_var);
      mul15_449 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_476_inst
    process(tmp13_427, tmp_415) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp13_427, tmp_415, tmp_var);
      tmp1_477 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_481_inst
    process(tmp1_477, tmp14_439) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_477, tmp14_439, tmp_var);
      tmp2_482 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_546_inst
    process(shl_535, conv27_542) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_535, conv27_542, tmp_var);
      add_547 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_564_inst
    process(shl29_553, conv32_560) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl29_553, conv32_560, tmp_var);
      add33_565 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_582_inst
    process(shl35_571, conv38_578) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl35_571, conv38_578, tmp_var);
      add39_583 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_600_inst
    process(shl41_589, conv44_596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl41_589, conv44_596, tmp_var);
      add45_601 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_618_inst
    process(shl47_607, conv50_614) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl47_607, conv50_614, tmp_var);
      add51_619 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_636_inst
    process(shl53_625, conv56_632) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl53_625, conv56_632, tmp_var);
      add57_637 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_654_inst
    process(shl59_643, conv62_650) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl59_643, conv62_650, tmp_var);
      add63_655 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_534_inst
    process(conv23_529) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv23_529, type_cast_533_wire_constant, tmp_var);
      shl_535 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_552_inst
    process(add_547) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_547, type_cast_551_wire_constant, tmp_var);
      shl29_553 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_570_inst
    process(add33_565) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add33_565, type_cast_569_wire_constant, tmp_var);
      shl35_571 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_588_inst
    process(add39_583) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add39_583, type_cast_587_wire_constant, tmp_var);
      shl41_589 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_606_inst
    process(add45_601) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add45_601, type_cast_605_wire_constant, tmp_var);
      shl47_607 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_624_inst
    process(add51_619) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add51_619, type_cast_623_wire_constant, tmp_var);
      shl53_625 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_642_inst
    process(add57_637) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add57_637, type_cast_641_wire_constant, tmp_var);
      shl59_643 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_497_inst
    process(tmp4_492) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp4_492, type_cast_496_wire_constant, tmp_var);
      tmp5_498 <= tmp_var; --
    end process;
    -- shared split operator group (24) : array_obj_ref_520_index_offset 
    ApIntAdd_group_24: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_519_scaled;
      array_obj_ref_520_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_520_index_offset_req_0;
      array_obj_ref_520_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_520_index_offset_req_1;
      array_obj_ref_520_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_24_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared load operator group (0) : ptr_deref_414_load_0 ptr_deref_426_load_0 ptr_deref_438_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_414_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_426_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_438_load_0_req_0;
      ptr_deref_414_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_426_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_438_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_414_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_426_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_438_load_0_req_1;
      ptr_deref_414_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_426_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_438_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_414_word_address_0 & ptr_deref_426_word_address_0 & ptr_deref_438_word_address_0;
      ptr_deref_414_data_0 <= data_out(95 downto 64);
      ptr_deref_426_data_0 <= data_out(63 downto 32);
      ptr_deref_438_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(6 downto 0),
          mtag => memory_space_5_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(31 downto 0),
          mtag => memory_space_5_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : STORE_col_high_332_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_col_high_332_store_0_req_0;
      STORE_col_high_332_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_col_high_332_store_0_req_1;
      STORE_col_high_332_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_col_high_332_word_address_0;
      data_in <= STORE_col_high_332_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(7 downto 0),
          mtag => memory_space_2_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : STORE_depth_high_338_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_depth_high_338_store_0_req_0;
      STORE_depth_high_338_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_depth_high_338_store_0_req_1;
      STORE_depth_high_338_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_depth_high_338_word_address_0;
      data_in <= STORE_depth_high_338_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(0 downto 0),
          mdata => memory_space_4_sr_data(7 downto 0),
          mtag => memory_space_4_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : STORE_pad_344_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_pad_344_store_0_req_0;
      STORE_pad_344_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_pad_344_store_0_req_1;
      STORE_pad_344_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_pad_344_word_address_0;
      data_in <= STORE_pad_344_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(7 downto 0),
          mtag => memory_space_7_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : STORE_row_high_326_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_row_high_326_store_0_req_0;
      STORE_row_high_326_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_row_high_326_store_0_req_1;
      STORE_row_high_326_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_row_high_326_word_address_0;
      data_in <= STORE_row_high_326_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(7 downto 0),
          mtag => memory_space_8_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_285_store_0 ptr_deref_303_store_0 ptr_deref_320_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_285_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_303_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_320_store_0_req_0;
      ptr_deref_285_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_303_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_320_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_285_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_303_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_320_store_0_req_1;
      ptr_deref_285_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_303_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_320_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup4_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_285_word_address_0 & ptr_deref_303_word_address_0 & ptr_deref_320_word_address_0;
      data_in <= ptr_deref_285_data_0 & ptr_deref_303_data_0 & ptr_deref_320_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(6 downto 0),
          mdata => memory_space_5_sr_data(31 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_363_store_0 ptr_deref_382_store_0 ptr_deref_401_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_363_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_382_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_401_store_0_req_0;
      ptr_deref_363_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_382_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_401_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_363_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_382_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_401_store_0_req_1;
      ptr_deref_363_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_382_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_401_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup5_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup5_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup5_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_363_word_address_0 & ptr_deref_382_word_address_0 & ptr_deref_401_word_address_0;
      data_in <= ptr_deref_363_data_0 & ptr_deref_382_data_0 & ptr_deref_401_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 3,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(6 downto 0),
          mdata => memory_space_6_sr_data(31 downto 0),
          mtag => memory_space_6_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_657_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_657_store_0_req_0;
      ptr_deref_657_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_657_store_0_req_1;
      ptr_deref_657_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_657_word_address_0;
      data_in <= ptr_deref_657_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared inport operator group (0) : RPIPE_zeropad_input_pipe_627_inst RPIPE_zeropad_input_pipe_645_inst RPIPE_zeropad_input_pipe_609_inst RPIPE_zeropad_input_pipe_591_inst RPIPE_zeropad_input_pipe_573_inst RPIPE_zeropad_input_pipe_290_inst RPIPE_zeropad_input_pipe_307_inst RPIPE_zeropad_input_pipe_324_inst RPIPE_zeropad_input_pipe_330_inst RPIPE_zeropad_input_pipe_336_inst RPIPE_zeropad_input_pipe_342_inst RPIPE_zeropad_input_pipe_348_inst RPIPE_zeropad_input_pipe_367_inst RPIPE_zeropad_input_pipe_386_inst RPIPE_zeropad_input_pipe_524_inst RPIPE_zeropad_input_pipe_537_inst RPIPE_zeropad_input_pipe_555_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(135 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 16 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 16 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 16 downto 0);
      signal guard_vector : std_logic_vector( 16 downto 0);
      constant outBUFs : IntegerArray(16 downto 0) := (16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(16 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false);
      constant guardBuffering: IntegerArray(16 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2);
      -- 
    begin -- 
      reqL_unguarded(16) <= RPIPE_zeropad_input_pipe_627_inst_req_0;
      reqL_unguarded(15) <= RPIPE_zeropad_input_pipe_645_inst_req_0;
      reqL_unguarded(14) <= RPIPE_zeropad_input_pipe_609_inst_req_0;
      reqL_unguarded(13) <= RPIPE_zeropad_input_pipe_591_inst_req_0;
      reqL_unguarded(12) <= RPIPE_zeropad_input_pipe_573_inst_req_0;
      reqL_unguarded(11) <= RPIPE_zeropad_input_pipe_290_inst_req_0;
      reqL_unguarded(10) <= RPIPE_zeropad_input_pipe_307_inst_req_0;
      reqL_unguarded(9) <= RPIPE_zeropad_input_pipe_324_inst_req_0;
      reqL_unguarded(8) <= RPIPE_zeropad_input_pipe_330_inst_req_0;
      reqL_unguarded(7) <= RPIPE_zeropad_input_pipe_336_inst_req_0;
      reqL_unguarded(6) <= RPIPE_zeropad_input_pipe_342_inst_req_0;
      reqL_unguarded(5) <= RPIPE_zeropad_input_pipe_348_inst_req_0;
      reqL_unguarded(4) <= RPIPE_zeropad_input_pipe_367_inst_req_0;
      reqL_unguarded(3) <= RPIPE_zeropad_input_pipe_386_inst_req_0;
      reqL_unguarded(2) <= RPIPE_zeropad_input_pipe_524_inst_req_0;
      reqL_unguarded(1) <= RPIPE_zeropad_input_pipe_537_inst_req_0;
      reqL_unguarded(0) <= RPIPE_zeropad_input_pipe_555_inst_req_0;
      RPIPE_zeropad_input_pipe_627_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_zeropad_input_pipe_645_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_zeropad_input_pipe_609_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_zeropad_input_pipe_591_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_zeropad_input_pipe_573_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_zeropad_input_pipe_290_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_zeropad_input_pipe_307_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_zeropad_input_pipe_324_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_zeropad_input_pipe_330_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_zeropad_input_pipe_336_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_zeropad_input_pipe_342_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_zeropad_input_pipe_348_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_zeropad_input_pipe_367_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_zeropad_input_pipe_386_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_zeropad_input_pipe_524_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_zeropad_input_pipe_537_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_zeropad_input_pipe_555_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(16) <= RPIPE_zeropad_input_pipe_627_inst_req_1;
      reqR_unguarded(15) <= RPIPE_zeropad_input_pipe_645_inst_req_1;
      reqR_unguarded(14) <= RPIPE_zeropad_input_pipe_609_inst_req_1;
      reqR_unguarded(13) <= RPIPE_zeropad_input_pipe_591_inst_req_1;
      reqR_unguarded(12) <= RPIPE_zeropad_input_pipe_573_inst_req_1;
      reqR_unguarded(11) <= RPIPE_zeropad_input_pipe_290_inst_req_1;
      reqR_unguarded(10) <= RPIPE_zeropad_input_pipe_307_inst_req_1;
      reqR_unguarded(9) <= RPIPE_zeropad_input_pipe_324_inst_req_1;
      reqR_unguarded(8) <= RPIPE_zeropad_input_pipe_330_inst_req_1;
      reqR_unguarded(7) <= RPIPE_zeropad_input_pipe_336_inst_req_1;
      reqR_unguarded(6) <= RPIPE_zeropad_input_pipe_342_inst_req_1;
      reqR_unguarded(5) <= RPIPE_zeropad_input_pipe_348_inst_req_1;
      reqR_unguarded(4) <= RPIPE_zeropad_input_pipe_367_inst_req_1;
      reqR_unguarded(3) <= RPIPE_zeropad_input_pipe_386_inst_req_1;
      reqR_unguarded(2) <= RPIPE_zeropad_input_pipe_524_inst_req_1;
      reqR_unguarded(1) <= RPIPE_zeropad_input_pipe_537_inst_req_1;
      reqR_unguarded(0) <= RPIPE_zeropad_input_pipe_555_inst_req_1;
      RPIPE_zeropad_input_pipe_627_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_zeropad_input_pipe_645_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_zeropad_input_pipe_609_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_zeropad_input_pipe_591_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_zeropad_input_pipe_573_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_zeropad_input_pipe_290_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_zeropad_input_pipe_307_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_zeropad_input_pipe_324_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_zeropad_input_pipe_330_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_zeropad_input_pipe_336_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_zeropad_input_pipe_342_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_zeropad_input_pipe_348_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_zeropad_input_pipe_367_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_zeropad_input_pipe_386_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_zeropad_input_pipe_524_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_zeropad_input_pipe_537_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_zeropad_input_pipe_555_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      call54_628 <= data_out(135 downto 128);
      call60_646 <= data_out(127 downto 120);
      call48_610 <= data_out(119 downto 112);
      call42_592 <= data_out(111 downto 104);
      call36_574 <= data_out(103 downto 96);
      call_291 <= data_out(95 downto 88);
      call1_308 <= data_out(87 downto 80);
      call3_325 <= data_out(79 downto 72);
      call4_331 <= data_out(71 downto 64);
      call5_337 <= data_out(63 downto 56);
      call6_343 <= data_out(55 downto 48);
      call7_349 <= data_out(47 downto 40);
      call9_368 <= data_out(39 downto 32);
      call11_387 <= data_out(31 downto 24);
      call22_525 <= data_out(23 downto 16);
      call25_538 <= data_out(15 downto 8);
      call30_556 <= data_out(7 downto 0);
      zeropad_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "zeropad_input_pipe_read_0_gI", nreqs => 17, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      zeropad_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "zeropad_input_pipe_read_0", data_width => 8,  num_reqs => 17,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => zeropad_input_pipe_pipe_read_req(0),
          oack => zeropad_input_pipe_pipe_read_ack(0),
          odata => zeropad_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(4 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_data : in   std_logic_vector(15 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D;
architecture zeropad3D_arch of zeropad3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_CP_2152_start: Boolean;
  signal zeropad3D_CP_2152_symbol: Boolean;
  -- volatile/operator module components. 
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(4 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(4 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_1026_inst_ack_1 : boolean;
  signal LOAD_row_high_941_load_0_req_0 : boolean;
  signal type_cast_975_inst_ack_1 : boolean;
  signal type_cast_975_inst_req_1 : boolean;
  signal LOAD_row_high_941_load_0_ack_0 : boolean;
  signal type_cast_975_inst_ack_0 : boolean;
  signal if_stmt_1016_branch_ack_1 : boolean;
  signal if_stmt_1016_branch_ack_0 : boolean;
  signal call_stmt_716_call_req_0 : boolean;
  signal call_stmt_716_call_ack_0 : boolean;
  signal call_stmt_716_call_req_1 : boolean;
  signal call_stmt_716_call_ack_1 : boolean;
  signal ptr_deref_727_load_0_req_0 : boolean;
  signal ptr_deref_727_load_0_ack_0 : boolean;
  signal ptr_deref_727_load_0_req_1 : boolean;
  signal ptr_deref_727_load_0_ack_1 : boolean;
  signal type_cast_731_inst_req_0 : boolean;
  signal type_cast_731_inst_ack_0 : boolean;
  signal type_cast_731_inst_req_1 : boolean;
  signal type_cast_731_inst_ack_1 : boolean;
  signal addr_of_1156_final_reg_ack_0 : boolean;
  signal if_stmt_1016_branch_req_0 : boolean;
  signal type_cast_1085_inst_ack_1 : boolean;
  signal type_cast_975_inst_req_0 : boolean;
  signal STORE_row_high_733_store_0_req_0 : boolean;
  signal STORE_row_high_733_store_0_ack_0 : boolean;
  signal STORE_row_high_733_store_0_req_1 : boolean;
  signal STORE_row_high_733_store_0_ack_1 : boolean;
  signal type_cast_996_inst_ack_1 : boolean;
  signal type_cast_1026_inst_req_1 : boolean;
  signal ptr_deref_746_load_0_req_0 : boolean;
  signal type_cast_996_inst_req_1 : boolean;
  signal ptr_deref_746_load_0_ack_0 : boolean;
  signal ptr_deref_746_load_0_req_1 : boolean;
  signal ptr_deref_746_load_0_ack_1 : boolean;
  signal type_cast_1085_inst_req_1 : boolean;
  signal addr_of_1156_final_reg_req_0 : boolean;
  signal type_cast_996_inst_ack_0 : boolean;
  signal type_cast_750_inst_req_0 : boolean;
  signal type_cast_750_inst_ack_0 : boolean;
  signal type_cast_1085_inst_ack_0 : boolean;
  signal type_cast_750_inst_req_1 : boolean;
  signal type_cast_750_inst_ack_1 : boolean;
  signal ptr_deref_1160_load_0_ack_0 : boolean;
  signal ptr_deref_1160_load_0_ack_1 : boolean;
  signal type_cast_996_inst_req_0 : boolean;
  signal type_cast_1085_inst_req_0 : boolean;
  signal type_cast_1066_inst_ack_1 : boolean;
  signal STORE_col_high_752_store_0_req_0 : boolean;
  signal STORE_col_high_752_store_0_ack_0 : boolean;
  signal STORE_col_high_752_store_0_req_1 : boolean;
  signal STORE_col_high_752_store_0_ack_1 : boolean;
  signal addr_of_1073_final_reg_ack_1 : boolean;
  signal LOAD_row_high_941_load_0_ack_1 : boolean;
  signal addr_of_1073_final_reg_req_1 : boolean;
  signal type_cast_1066_inst_req_1 : boolean;
  signal type_cast_1026_inst_ack_0 : boolean;
  signal if_stmt_965_branch_ack_0 : boolean;
  signal ptr_deref_765_load_0_req_0 : boolean;
  signal ptr_deref_765_load_0_ack_0 : boolean;
  signal type_cast_1026_inst_req_0 : boolean;
  signal ptr_deref_765_load_0_req_1 : boolean;
  signal ptr_deref_765_load_0_ack_1 : boolean;
  signal ptr_deref_1160_load_0_req_1 : boolean;
  signal LOAD_col_high_992_load_0_ack_1 : boolean;
  signal type_cast_1066_inst_ack_0 : boolean;
  signal type_cast_769_inst_req_0 : boolean;
  signal type_cast_1066_inst_req_0 : boolean;
  signal type_cast_769_inst_ack_0 : boolean;
  signal type_cast_769_inst_req_1 : boolean;
  signal type_cast_769_inst_ack_1 : boolean;
  signal ptr_deref_1160_load_0_req_0 : boolean;
  signal array_obj_ref_1155_index_offset_ack_1 : boolean;
  signal array_obj_ref_1155_index_offset_req_1 : boolean;
  signal addr_of_1073_final_reg_ack_0 : boolean;
  signal LOAD_col_high_992_load_0_req_1 : boolean;
  signal if_stmt_965_branch_ack_1 : boolean;
  signal STORE_depth_high_771_store_0_req_0 : boolean;
  signal STORE_depth_high_771_store_0_ack_0 : boolean;
  signal LOAD_row_high_941_load_0_req_1 : boolean;
  signal STORE_depth_high_771_store_0_req_1 : boolean;
  signal STORE_depth_high_771_store_0_ack_1 : boolean;
  signal addr_of_1073_final_reg_req_0 : boolean;
  signal type_cast_1149_inst_ack_1 : boolean;
  signal type_cast_1149_inst_req_1 : boolean;
  signal type_cast_1149_inst_ack_0 : boolean;
  signal array_obj_ref_1155_index_offset_ack_0 : boolean;
  signal addr_of_1156_final_reg_ack_1 : boolean;
  signal LOAD_pad_776_load_0_req_0 : boolean;
  signal LOAD_pad_776_load_0_ack_0 : boolean;
  signal if_stmt_965_branch_req_0 : boolean;
  signal addr_of_1156_final_reg_req_1 : boolean;
  signal LOAD_pad_776_load_0_req_1 : boolean;
  signal LOAD_pad_776_load_0_ack_1 : boolean;
  signal LOAD_col_high_992_load_0_ack_0 : boolean;
  signal array_obj_ref_1155_index_offset_req_0 : boolean;
  signal type_cast_1149_inst_req_0 : boolean;
  signal LOAD_col_high_992_load_0_req_0 : boolean;
  signal ptr_deref_1076_store_0_ack_1 : boolean;
  signal LOAD_depth_high_779_load_0_req_0 : boolean;
  signal LOAD_depth_high_779_load_0_ack_0 : boolean;
  signal LOAD_depth_high_779_load_0_req_1 : boolean;
  signal LOAD_depth_high_779_load_0_ack_1 : boolean;
  signal ptr_deref_1076_store_0_req_1 : boolean;
  signal LOAD_col_high_782_load_0_req_0 : boolean;
  signal LOAD_col_high_782_load_0_ack_0 : boolean;
  signal LOAD_col_high_782_load_0_req_1 : boolean;
  signal LOAD_col_high_782_load_0_ack_1 : boolean;
  signal array_obj_ref_1072_index_offset_ack_1 : boolean;
  signal array_obj_ref_1072_index_offset_req_1 : boolean;
  signal array_obj_ref_1072_index_offset_ack_0 : boolean;
  signal type_cast_1031_inst_ack_1 : boolean;
  signal type_cast_945_inst_ack_1 : boolean;
  signal type_cast_945_inst_req_1 : boolean;
  signal ptr_deref_794_load_0_req_0 : boolean;
  signal ptr_deref_794_load_0_ack_0 : boolean;
  signal ptr_deref_794_load_0_req_1 : boolean;
  signal if_stmt_984_branch_ack_0 : boolean;
  signal ptr_deref_794_load_0_ack_1 : boolean;
  signal array_obj_ref_1072_index_offset_req_0 : boolean;
  signal type_cast_1031_inst_req_1 : boolean;
  signal if_stmt_984_branch_ack_1 : boolean;
  signal type_cast_945_inst_ack_0 : boolean;
  signal type_cast_945_inst_req_0 : boolean;
  signal ptr_deref_806_load_0_req_0 : boolean;
  signal ptr_deref_806_load_0_ack_0 : boolean;
  signal ptr_deref_806_load_0_req_1 : boolean;
  signal ptr_deref_806_load_0_ack_1 : boolean;
  signal if_stmt_984_branch_req_0 : boolean;
  signal type_cast_1031_inst_ack_0 : boolean;
  signal type_cast_810_inst_req_0 : boolean;
  signal type_cast_1031_inst_req_0 : boolean;
  signal type_cast_810_inst_ack_0 : boolean;
  signal if_stmt_933_branch_ack_0 : boolean;
  signal type_cast_810_inst_req_1 : boolean;
  signal type_cast_810_inst_ack_1 : boolean;
  signal ptr_deref_1076_store_0_ack_0 : boolean;
  signal type_cast_814_inst_req_0 : boolean;
  signal type_cast_814_inst_ack_0 : boolean;
  signal ptr_deref_1076_store_0_req_0 : boolean;
  signal type_cast_814_inst_req_1 : boolean;
  signal type_cast_814_inst_ack_1 : boolean;
  signal type_cast_1560_inst_req_0 : boolean;
  signal type_cast_854_inst_req_0 : boolean;
  signal type_cast_854_inst_ack_0 : boolean;
  signal type_cast_854_inst_req_1 : boolean;
  signal type_cast_854_inst_ack_1 : boolean;
  signal type_cast_1560_inst_ack_0 : boolean;
  signal type_cast_924_inst_req_0 : boolean;
  signal type_cast_1706_inst_ack_0 : boolean;
  signal type_cast_924_inst_ack_0 : boolean;
  signal type_cast_924_inst_req_1 : boolean;
  signal type_cast_924_inst_ack_1 : boolean;
  signal if_stmt_933_branch_req_0 : boolean;
  signal if_stmt_933_branch_ack_1 : boolean;
  signal type_cast_1174_inst_req_0 : boolean;
  signal type_cast_1174_inst_ack_0 : boolean;
  signal type_cast_1174_inst_req_1 : boolean;
  signal type_cast_1174_inst_ack_1 : boolean;
  signal array_obj_ref_1180_index_offset_req_0 : boolean;
  signal array_obj_ref_1180_index_offset_ack_0 : boolean;
  signal array_obj_ref_1180_index_offset_req_1 : boolean;
  signal array_obj_ref_1180_index_offset_ack_1 : boolean;
  signal addr_of_1181_final_reg_req_0 : boolean;
  signal addr_of_1181_final_reg_ack_0 : boolean;
  signal addr_of_1181_final_reg_req_1 : boolean;
  signal addr_of_1181_final_reg_ack_1 : boolean;
  signal type_cast_1706_inst_req_0 : boolean;
  signal ptr_deref_1184_store_0_req_0 : boolean;
  signal ptr_deref_1184_store_0_ack_0 : boolean;
  signal ptr_deref_1184_store_0_req_1 : boolean;
  signal ptr_deref_1184_store_0_ack_1 : boolean;
  signal type_cast_1731_inst_ack_1 : boolean;
  signal type_cast_1192_inst_req_0 : boolean;
  signal type_cast_1192_inst_ack_0 : boolean;
  signal type_cast_1731_inst_req_1 : boolean;
  signal type_cast_1192_inst_req_1 : boolean;
  signal type_cast_1192_inst_ack_1 : boolean;
  signal LOAD_col_high_1556_load_0_ack_1 : boolean;
  signal if_stmt_1207_branch_req_0 : boolean;
  signal LOAD_col_high_1556_load_0_req_1 : boolean;
  signal if_stmt_1207_branch_ack_1 : boolean;
  signal if_stmt_1207_branch_ack_0 : boolean;
  signal addr_of_1713_final_reg_ack_0 : boolean;
  signal addr_of_1713_final_reg_req_0 : boolean;
  signal type_cast_1731_inst_ack_0 : boolean;
  signal type_cast_1231_inst_req_0 : boolean;
  signal type_cast_1231_inst_ack_0 : boolean;
  signal type_cast_1731_inst_req_0 : boolean;
  signal type_cast_1231_inst_req_1 : boolean;
  signal type_cast_1231_inst_ack_1 : boolean;
  signal type_cast_1642_inst_ack_1 : boolean;
  signal LOAD_col_high_1234_load_0_req_0 : boolean;
  signal LOAD_col_high_1234_load_0_ack_0 : boolean;
  signal LOAD_col_high_1556_load_0_ack_0 : boolean;
  signal LOAD_col_high_1556_load_0_req_0 : boolean;
  signal type_cast_1642_inst_req_1 : boolean;
  signal LOAD_col_high_1234_load_0_req_1 : boolean;
  signal LOAD_col_high_1234_load_0_ack_1 : boolean;
  signal ptr_deref_1741_store_0_ack_1 : boolean;
  signal if_stmt_1548_branch_ack_0 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal type_cast_1642_inst_ack_0 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal type_cast_1642_inst_req_0 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal array_obj_ref_1712_index_offset_ack_1 : boolean;
  signal type_cast_1258_inst_req_0 : boolean;
  signal type_cast_1258_inst_ack_0 : boolean;
  signal type_cast_1258_inst_req_1 : boolean;
  signal type_cast_1258_inst_ack_1 : boolean;
  signal ptr_deref_1741_store_0_ack_0 : boolean;
  signal addr_of_1738_final_reg_ack_1 : boolean;
  signal array_obj_ref_1712_index_offset_req_1 : boolean;
  signal type_cast_1275_inst_req_0 : boolean;
  signal type_cast_1275_inst_ack_0 : boolean;
  signal type_cast_1275_inst_req_1 : boolean;
  signal type_cast_1275_inst_ack_1 : boolean;
  signal addr_of_1738_final_reg_req_1 : boolean;
  signal ptr_deref_1741_store_0_req_0 : boolean;
  signal ptr_deref_1717_load_0_ack_1 : boolean;
  signal LOAD_row_high_1278_load_0_req_0 : boolean;
  signal LOAD_row_high_1278_load_0_ack_0 : boolean;
  signal if_stmt_1574_branch_ack_0 : boolean;
  signal LOAD_row_high_1278_load_0_req_1 : boolean;
  signal LOAD_row_high_1278_load_0_ack_1 : boolean;
  signal type_cast_1623_inst_ack_1 : boolean;
  signal ptr_deref_1741_store_0_req_1 : boolean;
  signal array_obj_ref_1712_index_offset_ack_0 : boolean;
  signal type_cast_1623_inst_req_1 : boolean;
  signal ptr_deref_1717_load_0_req_1 : boolean;
  signal type_cast_1282_inst_req_0 : boolean;
  signal type_cast_1282_inst_ack_0 : boolean;
  signal type_cast_1282_inst_req_1 : boolean;
  signal ptr_deref_1633_store_0_ack_1 : boolean;
  signal type_cast_1282_inst_ack_1 : boolean;
  signal addr_of_1738_final_reg_ack_0 : boolean;
  signal ptr_deref_1633_store_0_req_1 : boolean;
  signal if_stmt_1300_branch_req_0 : boolean;
  signal if_stmt_1300_branch_ack_1 : boolean;
  signal addr_of_1630_final_reg_ack_1 : boolean;
  signal if_stmt_1300_branch_ack_0 : boolean;
  signal addr_of_1630_final_reg_req_1 : boolean;
  signal array_obj_ref_1712_index_offset_req_0 : boolean;
  signal type_cast_1340_inst_req_0 : boolean;
  signal type_cast_1340_inst_ack_0 : boolean;
  signal type_cast_1340_inst_req_1 : boolean;
  signal type_cast_1340_inst_ack_1 : boolean;
  signal addr_of_1738_final_reg_req_0 : boolean;
  signal type_cast_1623_inst_ack_0 : boolean;
  signal ptr_deref_1717_load_0_ack_0 : boolean;
  signal ptr_deref_1717_load_0_req_0 : boolean;
  signal LOAD_pad_1349_load_0_req_0 : boolean;
  signal type_cast_1623_inst_req_0 : boolean;
  signal LOAD_pad_1349_load_0_ack_0 : boolean;
  signal if_stmt_1574_branch_ack_1 : boolean;
  signal LOAD_pad_1349_load_0_req_1 : boolean;
  signal LOAD_pad_1349_load_0_ack_1 : boolean;
  signal LOAD_depth_high_1352_load_0_req_0 : boolean;
  signal LOAD_depth_high_1352_load_0_ack_0 : boolean;
  signal LOAD_depth_high_1352_load_0_req_1 : boolean;
  signal type_cast_1589_inst_ack_1 : boolean;
  signal LOAD_depth_high_1352_load_0_ack_1 : boolean;
  signal addr_of_1630_final_reg_ack_0 : boolean;
  signal type_cast_1589_inst_req_1 : boolean;
  signal type_cast_1589_inst_ack_0 : boolean;
  signal addr_of_1630_final_reg_req_0 : boolean;
  signal ptr_deref_1633_store_0_ack_0 : boolean;
  signal if_stmt_1574_branch_req_0 : boolean;
  signal ptr_deref_1364_load_0_req_0 : boolean;
  signal type_cast_1589_inst_req_0 : boolean;
  signal ptr_deref_1364_load_0_ack_0 : boolean;
  signal ptr_deref_1364_load_0_req_1 : boolean;
  signal ptr_deref_1364_load_0_ack_1 : boolean;
  signal array_obj_ref_1737_index_offset_ack_1 : boolean;
  signal array_obj_ref_1737_index_offset_req_1 : boolean;
  signal ptr_deref_1633_store_0_req_0 : boolean;
  signal ptr_deref_1376_load_0_req_0 : boolean;
  signal ptr_deref_1376_load_0_ack_0 : boolean;
  signal type_cast_1560_inst_ack_1 : boolean;
  signal ptr_deref_1376_load_0_req_1 : boolean;
  signal type_cast_1584_inst_ack_1 : boolean;
  signal ptr_deref_1376_load_0_ack_1 : boolean;
  signal type_cast_1584_inst_req_1 : boolean;
  signal if_stmt_1548_branch_ack_1 : boolean;
  signal type_cast_1380_inst_req_0 : boolean;
  signal type_cast_1380_inst_ack_0 : boolean;
  signal type_cast_1380_inst_req_1 : boolean;
  signal type_cast_1380_inst_ack_1 : boolean;
  signal array_obj_ref_1737_index_offset_ack_0 : boolean;
  signal array_obj_ref_1737_index_offset_req_0 : boolean;
  signal type_cast_1706_inst_ack_1 : boolean;
  signal type_cast_1419_inst_req_0 : boolean;
  signal type_cast_1419_inst_ack_0 : boolean;
  signal type_cast_1419_inst_req_1 : boolean;
  signal type_cast_1419_inst_ack_1 : boolean;
  signal type_cast_1584_inst_ack_0 : boolean;
  signal type_cast_1706_inst_req_1 : boolean;
  signal type_cast_1488_inst_req_0 : boolean;
  signal type_cast_1488_inst_ack_0 : boolean;
  signal type_cast_1488_inst_req_1 : boolean;
  signal type_cast_1488_inst_ack_1 : boolean;
  signal type_cast_1584_inst_req_0 : boolean;
  signal array_obj_ref_1629_index_offset_ack_1 : boolean;
  signal if_stmt_1497_branch_req_0 : boolean;
  signal array_obj_ref_1629_index_offset_req_1 : boolean;
  signal if_stmt_1497_branch_ack_1 : boolean;
  signal if_stmt_1497_branch_ack_0 : boolean;
  signal addr_of_1713_final_reg_ack_1 : boolean;
  signal type_cast_1560_inst_req_1 : boolean;
  signal array_obj_ref_1629_index_offset_ack_0 : boolean;
  signal addr_of_1713_final_reg_req_1 : boolean;
  signal LOAD_row_high_1505_load_0_req_0 : boolean;
  signal LOAD_row_high_1505_load_0_ack_0 : boolean;
  signal LOAD_row_high_1505_load_0_req_1 : boolean;
  signal LOAD_row_high_1505_load_0_ack_1 : boolean;
  signal array_obj_ref_1629_index_offset_req_0 : boolean;
  signal type_cast_1509_inst_req_0 : boolean;
  signal type_cast_1509_inst_ack_0 : boolean;
  signal type_cast_1509_inst_req_1 : boolean;
  signal type_cast_1509_inst_ack_1 : boolean;
  signal ptr_deref_2189_store_0_req_1 : boolean;
  signal if_stmt_1529_branch_req_0 : boolean;
  signal if_stmt_1529_branch_ack_1 : boolean;
  signal if_stmt_1529_branch_ack_0 : boolean;
  signal ptr_deref_2189_store_0_ack_1 : boolean;
  signal type_cast_1539_inst_req_0 : boolean;
  signal type_cast_1539_inst_ack_0 : boolean;
  signal type_cast_1539_inst_req_1 : boolean;
  signal type_cast_1539_inst_ack_1 : boolean;
  signal if_stmt_1548_branch_req_0 : boolean;
  signal type_cast_3012_inst_req_0 : boolean;
  signal type_cast_3012_inst_ack_0 : boolean;
  signal type_cast_3012_inst_req_1 : boolean;
  signal type_cast_3012_inst_ack_1 : boolean;
  signal phi_stmt_3009_req_0 : boolean;
  signal phi_stmt_3005_ack_0 : boolean;
  signal phi_stmt_3009_ack_0 : boolean;
  signal type_cast_1749_inst_req_0 : boolean;
  signal type_cast_1749_inst_ack_0 : boolean;
  signal type_cast_1749_inst_req_1 : boolean;
  signal type_cast_1749_inst_ack_1 : boolean;
  signal if_stmt_1764_branch_req_0 : boolean;
  signal if_stmt_1764_branch_ack_1 : boolean;
  signal if_stmt_1764_branch_ack_0 : boolean;
  signal type_cast_1788_inst_req_0 : boolean;
  signal type_cast_1788_inst_ack_0 : boolean;
  signal type_cast_1788_inst_req_1 : boolean;
  signal type_cast_1788_inst_ack_1 : boolean;
  signal type_cast_2198_inst_ack_1 : boolean;
  signal LOAD_col_high_1791_load_0_req_0 : boolean;
  signal LOAD_col_high_1791_load_0_ack_0 : boolean;
  signal type_cast_2198_inst_req_1 : boolean;
  signal LOAD_col_high_1791_load_0_req_1 : boolean;
  signal LOAD_col_high_1791_load_0_ack_1 : boolean;
  signal type_cast_2198_inst_ack_0 : boolean;
  signal type_cast_2198_inst_req_0 : boolean;
  signal ptr_deref_2297_store_0_ack_1 : boolean;
  signal type_cast_2344_inst_ack_0 : boolean;
  signal type_cast_1795_inst_req_0 : boolean;
  signal type_cast_1795_inst_ack_0 : boolean;
  signal type_cast_2344_inst_req_0 : boolean;
  signal type_cast_1795_inst_req_1 : boolean;
  signal type_cast_1795_inst_ack_1 : boolean;
  signal ptr_deref_2297_store_0_req_1 : boolean;
  signal type_cast_1809_inst_req_0 : boolean;
  signal type_cast_1809_inst_ack_0 : boolean;
  signal type_cast_1809_inst_req_1 : boolean;
  signal addr_of_2294_final_reg_ack_1 : boolean;
  signal type_cast_1809_inst_ack_1 : boolean;
  signal LOAD_col_high_2347_load_0_ack_0 : boolean;
  signal LOAD_col_high_2347_load_0_req_0 : boolean;
  signal addr_of_2294_final_reg_req_1 : boolean;
  signal type_cast_1825_inst_req_0 : boolean;
  signal type_cast_1825_inst_ack_0 : boolean;
  signal type_cast_1825_inst_req_1 : boolean;
  signal type_cast_1825_inst_ack_1 : boolean;
  signal ptr_deref_2273_load_0_ack_1 : boolean;
  signal ptr_deref_2273_load_0_req_1 : boolean;
  signal LOAD_row_high_1828_load_0_req_0 : boolean;
  signal LOAD_row_high_1828_load_0_ack_0 : boolean;
  signal LOAD_row_high_1828_load_0_req_1 : boolean;
  signal LOAD_row_high_1828_load_0_ack_1 : boolean;
  signal LOAD_col_high_2347_load_0_ack_1 : boolean;
  signal ptr_deref_2297_store_0_ack_0 : boolean;
  signal addr_of_2294_final_reg_ack_0 : boolean;
  signal type_cast_1832_inst_req_0 : boolean;
  signal addr_of_2294_final_reg_req_0 : boolean;
  signal type_cast_1832_inst_ack_0 : boolean;
  signal if_stmt_2320_branch_ack_0 : boolean;
  signal type_cast_1832_inst_req_1 : boolean;
  signal type_cast_1832_inst_ack_1 : boolean;
  signal if_stmt_1850_branch_req_0 : boolean;
  signal if_stmt_1850_branch_ack_1 : boolean;
  signal if_stmt_1850_branch_ack_0 : boolean;
  signal type_cast_2287_inst_ack_1 : boolean;
  signal type_cast_2287_inst_req_1 : boolean;
  signal ptr_deref_2297_store_0_req_0 : boolean;
  signal type_cast_1890_inst_req_0 : boolean;
  signal type_cast_1890_inst_ack_0 : boolean;
  signal if_stmt_2320_branch_ack_1 : boolean;
  signal type_cast_1890_inst_req_1 : boolean;
  signal type_cast_1890_inst_ack_1 : boolean;
  signal type_cast_2344_inst_ack_1 : boolean;
  signal ptr_deref_2273_load_0_ack_0 : boolean;
  signal LOAD_pad_1899_load_0_req_0 : boolean;
  signal ptr_deref_2273_load_0_req_0 : boolean;
  signal LOAD_pad_1899_load_0_ack_0 : boolean;
  signal LOAD_pad_1899_load_0_req_1 : boolean;
  signal LOAD_pad_1899_load_0_ack_1 : boolean;
  signal if_stmt_2320_branch_req_0 : boolean;
  signal LOAD_col_high_2347_load_0_req_1 : boolean;
  signal LOAD_depth_high_1902_load_0_req_0 : boolean;
  signal LOAD_depth_high_1902_load_0_ack_0 : boolean;
  signal LOAD_depth_high_1902_load_0_req_1 : boolean;
  signal LOAD_depth_high_1902_load_0_ack_1 : boolean;
  signal type_cast_2344_inst_req_1 : boolean;
  signal array_obj_ref_2293_index_offset_ack_1 : boolean;
  signal array_obj_ref_2293_index_offset_req_1 : boolean;
  signal type_cast_2287_inst_ack_0 : boolean;
  signal ptr_deref_1914_load_0_req_0 : boolean;
  signal ptr_deref_1914_load_0_ack_0 : boolean;
  signal ptr_deref_1914_load_0_req_1 : boolean;
  signal ptr_deref_1914_load_0_ack_1 : boolean;
  signal array_obj_ref_2293_index_offset_ack_0 : boolean;
  signal array_obj_ref_2293_index_offset_req_0 : boolean;
  signal ptr_deref_2189_store_0_ack_0 : boolean;
  signal addr_of_2269_final_reg_ack_1 : boolean;
  signal ptr_deref_1926_load_0_req_0 : boolean;
  signal addr_of_2269_final_reg_req_1 : boolean;
  signal ptr_deref_1926_load_0_ack_0 : boolean;
  signal ptr_deref_2189_store_0_req_0 : boolean;
  signal ptr_deref_1926_load_0_req_1 : boolean;
  signal ptr_deref_1926_load_0_ack_1 : boolean;
  signal type_cast_2262_inst_ack_1 : boolean;
  signal addr_of_2269_final_reg_ack_0 : boolean;
  signal addr_of_2269_final_reg_req_0 : boolean;
  signal type_cast_1930_inst_req_0 : boolean;
  signal type_cast_1930_inst_ack_0 : boolean;
  signal type_cast_1930_inst_req_1 : boolean;
  signal type_cast_1930_inst_ack_1 : boolean;
  signal type_cast_2262_inst_req_1 : boolean;
  signal type_cast_2305_inst_ack_1 : boolean;
  signal type_cast_1969_inst_req_0 : boolean;
  signal type_cast_1969_inst_ack_0 : boolean;
  signal type_cast_2305_inst_req_1 : boolean;
  signal type_cast_1969_inst_req_1 : boolean;
  signal type_cast_1969_inst_ack_1 : boolean;
  signal type_cast_2262_inst_ack_0 : boolean;
  signal type_cast_2038_inst_req_0 : boolean;
  signal type_cast_2038_inst_ack_0 : boolean;
  signal type_cast_2038_inst_req_1 : boolean;
  signal type_cast_2038_inst_ack_1 : boolean;
  signal type_cast_2262_inst_req_0 : boolean;
  signal array_obj_ref_2268_index_offset_ack_1 : boolean;
  signal type_cast_2305_inst_ack_0 : boolean;
  signal type_cast_2287_inst_req_0 : boolean;
  signal type_cast_2305_inst_req_0 : boolean;
  signal if_stmt_2047_branch_req_0 : boolean;
  signal array_obj_ref_2268_index_offset_req_1 : boolean;
  signal if_stmt_2047_branch_ack_1 : boolean;
  signal if_stmt_2047_branch_ack_0 : boolean;
  signal array_obj_ref_2268_index_offset_ack_0 : boolean;
  signal LOAD_row_high_2055_load_0_req_0 : boolean;
  signal array_obj_ref_2268_index_offset_req_0 : boolean;
  signal LOAD_row_high_2055_load_0_ack_0 : boolean;
  signal LOAD_row_high_2055_load_0_req_1 : boolean;
  signal LOAD_row_high_2055_load_0_ack_1 : boolean;
  signal type_cast_2059_inst_req_0 : boolean;
  signal type_cast_2059_inst_ack_0 : boolean;
  signal LOAD_row_high_2954_load_0_req_0 : boolean;
  signal type_cast_2059_inst_req_1 : boolean;
  signal type_cast_2059_inst_ack_1 : boolean;
  signal addr_of_2864_final_reg_req_0 : boolean;
  signal if_stmt_2079_branch_req_0 : boolean;
  signal if_stmt_2079_branch_ack_1 : boolean;
  signal if_stmt_2079_branch_ack_0 : boolean;
  signal type_cast_2921_inst_req_1 : boolean;
  signal type_cast_2089_inst_req_0 : boolean;
  signal type_cast_2089_inst_ack_0 : boolean;
  signal type_cast_2089_inst_req_1 : boolean;
  signal type_cast_2914_inst_req_0 : boolean;
  signal type_cast_2089_inst_ack_1 : boolean;
  signal type_cast_2921_inst_ack_1 : boolean;
  signal type_cast_2857_inst_req_0 : boolean;
  signal if_stmt_2098_branch_req_0 : boolean;
  signal if_stmt_2098_branch_ack_1 : boolean;
  signal if_stmt_2098_branch_ack_0 : boolean;
  signal type_cast_2914_inst_ack_0 : boolean;
  signal LOAD_col_high_2106_load_0_req_0 : boolean;
  signal LOAD_col_high_2106_load_0_ack_0 : boolean;
  signal LOAD_col_high_2106_load_0_req_1 : boolean;
  signal type_cast_2914_inst_req_1 : boolean;
  signal LOAD_col_high_2106_load_0_ack_1 : boolean;
  signal addr_of_2864_final_reg_ack_0 : boolean;
  signal type_cast_2110_inst_req_0 : boolean;
  signal type_cast_2110_inst_ack_0 : boolean;
  signal type_cast_2110_inst_req_1 : boolean;
  signal type_cast_2110_inst_ack_1 : boolean;
  signal type_cast_2914_inst_ack_1 : boolean;
  signal type_cast_2857_inst_ack_0 : boolean;
  signal if_stmt_2130_branch_req_0 : boolean;
  signal if_stmt_2130_branch_ack_1 : boolean;
  signal if_stmt_2130_branch_ack_0 : boolean;
  signal type_cast_2140_inst_req_0 : boolean;
  signal type_cast_2140_inst_ack_0 : boolean;
  signal type_cast_2140_inst_req_1 : boolean;
  signal type_cast_2140_inst_ack_1 : boolean;
  signal type_cast_2145_inst_req_0 : boolean;
  signal type_cast_2145_inst_ack_0 : boolean;
  signal type_cast_2145_inst_req_1 : boolean;
  signal type_cast_2145_inst_ack_1 : boolean;
  signal type_cast_2179_inst_req_0 : boolean;
  signal type_cast_2179_inst_ack_0 : boolean;
  signal type_cast_2179_inst_req_1 : boolean;
  signal type_cast_2179_inst_ack_1 : boolean;
  signal array_obj_ref_2185_index_offset_req_0 : boolean;
  signal array_obj_ref_2185_index_offset_ack_0 : boolean;
  signal array_obj_ref_2185_index_offset_req_1 : boolean;
  signal array_obj_ref_2185_index_offset_ack_1 : boolean;
  signal addr_of_2186_final_reg_req_0 : boolean;
  signal addr_of_2186_final_reg_ack_0 : boolean;
  signal addr_of_2186_final_reg_req_1 : boolean;
  signal addr_of_2186_final_reg_ack_1 : boolean;
  signal type_cast_2351_inst_req_0 : boolean;
  signal type_cast_2351_inst_ack_0 : boolean;
  signal type_cast_2351_inst_req_1 : boolean;
  signal type_cast_2351_inst_ack_1 : boolean;
  signal type_cast_2371_inst_req_0 : boolean;
  signal type_cast_2371_inst_ack_0 : boolean;
  signal type_cast_2371_inst_req_1 : boolean;
  signal type_cast_2371_inst_ack_1 : boolean;
  signal type_cast_2388_inst_req_0 : boolean;
  signal type_cast_2388_inst_ack_0 : boolean;
  signal type_cast_2388_inst_req_1 : boolean;
  signal type_cast_2388_inst_ack_1 : boolean;
  signal LOAD_row_high_2391_load_0_req_0 : boolean;
  signal LOAD_row_high_2391_load_0_ack_0 : boolean;
  signal LOAD_row_high_2391_load_0_req_1 : boolean;
  signal LOAD_row_high_2391_load_0_ack_1 : boolean;
  signal type_cast_2395_inst_req_0 : boolean;
  signal type_cast_2395_inst_ack_0 : boolean;
  signal type_cast_2395_inst_req_1 : boolean;
  signal type_cast_2395_inst_ack_1 : boolean;
  signal if_stmt_2413_branch_req_0 : boolean;
  signal if_stmt_2413_branch_ack_1 : boolean;
  signal if_stmt_2413_branch_ack_0 : boolean;
  signal type_cast_2457_inst_req_0 : boolean;
  signal type_cast_2457_inst_ack_0 : boolean;
  signal type_cast_2457_inst_req_1 : boolean;
  signal type_cast_2457_inst_ack_1 : boolean;
  signal type_cast_2467_inst_req_0 : boolean;
  signal type_cast_2467_inst_ack_0 : boolean;
  signal type_cast_2467_inst_req_1 : boolean;
  signal type_cast_2467_inst_ack_1 : boolean;
  signal LOAD_row_high_2954_load_0_ack_1 : boolean;
  signal type_cast_2935_inst_ack_1 : boolean;
  signal type_cast_2935_inst_req_1 : boolean;
  signal LOAD_pad_2476_load_0_req_0 : boolean;
  signal LOAD_pad_2476_load_0_ack_0 : boolean;
  signal LOAD_pad_2476_load_0_req_1 : boolean;
  signal LOAD_pad_2476_load_0_ack_1 : boolean;
  signal LOAD_row_high_2954_load_0_req_1 : boolean;
  signal if_stmt_2890_branch_ack_0 : boolean;
  signal if_stmt_2890_branch_ack_1 : boolean;
  signal LOAD_depth_high_2479_load_0_req_0 : boolean;
  signal LOAD_depth_high_2479_load_0_ack_0 : boolean;
  signal if_stmt_2890_branch_req_0 : boolean;
  signal LOAD_depth_high_2479_load_0_req_1 : boolean;
  signal LOAD_depth_high_2479_load_0_ack_1 : boolean;
  signal type_cast_2875_inst_ack_1 : boolean;
  signal type_cast_2875_inst_req_1 : boolean;
  signal type_cast_2921_inst_ack_0 : boolean;
  signal type_cast_2921_inst_req_0 : boolean;
  signal ptr_deref_2491_load_0_req_0 : boolean;
  signal type_cast_2875_inst_ack_0 : boolean;
  signal ptr_deref_2491_load_0_ack_0 : boolean;
  signal ptr_deref_2491_load_0_req_1 : boolean;
  signal type_cast_2875_inst_req_0 : boolean;
  signal ptr_deref_2491_load_0_ack_1 : boolean;
  signal ptr_deref_2867_store_0_ack_1 : boolean;
  signal ptr_deref_2867_store_0_req_1 : boolean;
  signal addr_of_2864_final_reg_ack_1 : boolean;
  signal ptr_deref_2503_load_0_req_0 : boolean;
  signal ptr_deref_2503_load_0_ack_0 : boolean;
  signal ptr_deref_2843_load_0_ack_1 : boolean;
  signal addr_of_2864_final_reg_req_1 : boolean;
  signal ptr_deref_2503_load_0_req_1 : boolean;
  signal ptr_deref_2503_load_0_ack_1 : boolean;
  signal array_obj_ref_2863_index_offset_ack_1 : boolean;
  signal type_cast_2935_inst_ack_0 : boolean;
  signal array_obj_ref_2863_index_offset_req_1 : boolean;
  signal ptr_deref_2843_load_0_req_1 : boolean;
  signal type_cast_2951_inst_ack_0 : boolean;
  signal ptr_deref_2867_store_0_ack_0 : boolean;
  signal ptr_deref_2867_store_0_req_0 : boolean;
  signal type_cast_2507_inst_req_0 : boolean;
  signal type_cast_2507_inst_ack_0 : boolean;
  signal type_cast_2507_inst_req_1 : boolean;
  signal type_cast_2507_inst_ack_1 : boolean;
  signal type_cast_2935_inst_req_0 : boolean;
  signal LOAD_col_high_2917_load_0_ack_1 : boolean;
  signal type_cast_2546_inst_req_0 : boolean;
  signal LOAD_col_high_2917_load_0_req_1 : boolean;
  signal type_cast_2546_inst_ack_0 : boolean;
  signal type_cast_2546_inst_req_1 : boolean;
  signal type_cast_2546_inst_ack_1 : boolean;
  signal type_cast_2857_inst_ack_1 : boolean;
  signal type_cast_2857_inst_req_1 : boolean;
  signal type_cast_2614_inst_req_0 : boolean;
  signal type_cast_2614_inst_ack_0 : boolean;
  signal type_cast_2614_inst_req_1 : boolean;
  signal type_cast_2614_inst_ack_1 : boolean;
  signal array_obj_ref_2863_index_offset_ack_0 : boolean;
  signal array_obj_ref_2863_index_offset_req_0 : boolean;
  signal type_cast_2951_inst_req_0 : boolean;
  signal if_stmt_2623_branch_req_0 : boolean;
  signal if_stmt_2623_branch_ack_1 : boolean;
  signal if_stmt_2623_branch_ack_0 : boolean;
  signal LOAD_row_high_2631_load_0_req_0 : boolean;
  signal LOAD_row_high_2631_load_0_ack_0 : boolean;
  signal LOAD_row_high_2631_load_0_req_1 : boolean;
  signal LOAD_row_high_2631_load_0_ack_1 : boolean;
  signal LOAD_row_high_2954_load_0_ack_0 : boolean;
  signal type_cast_2635_inst_req_0 : boolean;
  signal LOAD_col_high_2917_load_0_ack_0 : boolean;
  signal type_cast_2635_inst_ack_0 : boolean;
  signal type_cast_2951_inst_ack_1 : boolean;
  signal type_cast_2635_inst_req_1 : boolean;
  signal LOAD_col_high_2917_load_0_req_0 : boolean;
  signal type_cast_2635_inst_ack_1 : boolean;
  signal if_stmt_2655_branch_req_0 : boolean;
  signal if_stmt_2655_branch_ack_1 : boolean;
  signal ptr_deref_3429_store_0_req_0 : boolean;
  signal if_stmt_2655_branch_ack_0 : boolean;
  signal type_cast_3503_inst_req_0 : boolean;
  signal type_cast_3503_inst_ack_0 : boolean;
  signal type_cast_3595_inst_req_0 : boolean;
  signal type_cast_2665_inst_req_0 : boolean;
  signal type_cast_2665_inst_ack_0 : boolean;
  signal type_cast_3595_inst_ack_0 : boolean;
  signal type_cast_2665_inst_req_1 : boolean;
  signal type_cast_2665_inst_ack_1 : boolean;
  signal ptr_deref_3429_store_0_ack_0 : boolean;
  signal type_cast_3503_inst_req_1 : boolean;
  signal if_stmt_2674_branch_req_0 : boolean;
  signal if_stmt_2674_branch_ack_1 : boolean;
  signal if_stmt_2674_branch_ack_0 : boolean;
  signal LOAD_col_high_2682_load_0_req_0 : boolean;
  signal LOAD_col_high_2682_load_0_ack_0 : boolean;
  signal LOAD_col_high_2682_load_0_req_1 : boolean;
  signal LOAD_col_high_2682_load_0_ack_1 : boolean;
  signal type_cast_3527_inst_req_1 : boolean;
  signal LOAD_col_high_3479_load_0_req_1 : boolean;
  signal type_cast_2686_inst_req_0 : boolean;
  signal type_cast_2686_inst_ack_0 : boolean;
  signal type_cast_2686_inst_req_1 : boolean;
  signal LOAD_col_high_3479_load_0_ack_1 : boolean;
  signal type_cast_2686_inst_ack_1 : boolean;
  signal type_cast_3595_inst_req_1 : boolean;
  signal type_cast_3437_inst_req_0 : boolean;
  signal if_stmt_2700_branch_req_0 : boolean;
  signal type_cast_3503_inst_ack_1 : boolean;
  signal if_stmt_2700_branch_ack_1 : boolean;
  signal if_stmt_2700_branch_ack_0 : boolean;
  signal type_cast_2710_inst_req_0 : boolean;
  signal type_cast_2710_inst_ack_0 : boolean;
  signal type_cast_3595_inst_ack_1 : boolean;
  signal type_cast_2710_inst_req_1 : boolean;
  signal type_cast_2710_inst_ack_1 : boolean;
  signal type_cast_3437_inst_ack_0 : boolean;
  signal type_cast_2715_inst_req_0 : boolean;
  signal type_cast_2715_inst_ack_0 : boolean;
  signal type_cast_2715_inst_req_1 : boolean;
  signal type_cast_2715_inst_ack_1 : boolean;
  signal type_cast_2749_inst_req_0 : boolean;
  signal type_cast_2749_inst_ack_0 : boolean;
  signal type_cast_2749_inst_req_1 : boolean;
  signal type_cast_2749_inst_ack_1 : boolean;
  signal if_stmt_3452_branch_req_0 : boolean;
  signal type_cast_3527_inst_ack_1 : boolean;
  signal array_obj_ref_2755_index_offset_req_0 : boolean;
  signal array_obj_ref_2755_index_offset_ack_0 : boolean;
  signal array_obj_ref_2755_index_offset_req_1 : boolean;
  signal array_obj_ref_2755_index_offset_ack_1 : boolean;
  signal addr_of_2756_final_reg_req_0 : boolean;
  signal addr_of_2756_final_reg_ack_0 : boolean;
  signal addr_of_2756_final_reg_req_1 : boolean;
  signal addr_of_2756_final_reg_ack_1 : boolean;
  signal ptr_deref_2759_store_0_req_0 : boolean;
  signal ptr_deref_2759_store_0_ack_0 : boolean;
  signal ptr_deref_2759_store_0_req_1 : boolean;
  signal ptr_deref_2759_store_0_ack_1 : boolean;
  signal type_cast_2768_inst_req_0 : boolean;
  signal type_cast_2768_inst_ack_0 : boolean;
  signal type_cast_2768_inst_req_1 : boolean;
  signal type_cast_2768_inst_ack_1 : boolean;
  signal type_cast_2832_inst_req_0 : boolean;
  signal type_cast_2832_inst_ack_0 : boolean;
  signal type_cast_2832_inst_req_1 : boolean;
  signal type_cast_2832_inst_ack_1 : boolean;
  signal array_obj_ref_2838_index_offset_req_0 : boolean;
  signal array_obj_ref_2838_index_offset_ack_0 : boolean;
  signal array_obj_ref_2838_index_offset_req_1 : boolean;
  signal array_obj_ref_2838_index_offset_ack_1 : boolean;
  signal addr_of_2839_final_reg_req_0 : boolean;
  signal addr_of_2839_final_reg_ack_0 : boolean;
  signal addr_of_2839_final_reg_req_1 : boolean;
  signal addr_of_2839_final_reg_ack_1 : boolean;
  signal type_cast_2951_inst_req_1 : boolean;
  signal ptr_deref_2843_load_0_req_0 : boolean;
  signal ptr_deref_2843_load_0_ack_0 : boolean;
  signal type_cast_2958_inst_req_0 : boolean;
  signal type_cast_2958_inst_ack_0 : boolean;
  signal type_cast_2958_inst_req_1 : boolean;
  signal type_cast_2958_inst_ack_1 : boolean;
  signal if_stmt_2976_branch_req_0 : boolean;
  signal if_stmt_2976_branch_ack_1 : boolean;
  signal if_stmt_2976_branch_ack_0 : boolean;
  signal type_cast_3016_inst_req_0 : boolean;
  signal type_cast_3016_inst_ack_0 : boolean;
  signal type_cast_3016_inst_req_1 : boolean;
  signal type_cast_3016_inst_ack_1 : boolean;
  signal LOAD_pad_3025_load_0_req_0 : boolean;
  signal LOAD_pad_3025_load_0_ack_0 : boolean;
  signal LOAD_pad_3025_load_0_req_1 : boolean;
  signal LOAD_pad_3025_load_0_ack_1 : boolean;
  signal LOAD_depth_high_3028_load_0_req_0 : boolean;
  signal LOAD_depth_high_3028_load_0_ack_0 : boolean;
  signal LOAD_depth_high_3028_load_0_req_1 : boolean;
  signal LOAD_depth_high_3028_load_0_ack_1 : boolean;
  signal ptr_deref_3040_load_0_req_0 : boolean;
  signal ptr_deref_3040_load_0_ack_0 : boolean;
  signal ptr_deref_3040_load_0_req_1 : boolean;
  signal ptr_deref_3040_load_0_ack_1 : boolean;
  signal ptr_deref_3052_load_0_req_0 : boolean;
  signal ptr_deref_3052_load_0_ack_0 : boolean;
  signal ptr_deref_3052_load_0_req_1 : boolean;
  signal ptr_deref_3052_load_0_ack_1 : boolean;
  signal LOAD_col_high_3479_load_0_ack_0 : boolean;
  signal LOAD_col_high_3479_load_0_req_0 : boolean;
  signal type_cast_3056_inst_req_0 : boolean;
  signal LOAD_row_high_3523_load_0_ack_0 : boolean;
  signal type_cast_3056_inst_ack_0 : boolean;
  signal type_cast_3056_inst_req_1 : boolean;
  signal LOAD_row_high_3523_load_0_req_0 : boolean;
  signal type_cast_3056_inst_ack_1 : boolean;
  signal type_cast_3605_inst_ack_1 : boolean;
  signal type_cast_3605_inst_req_1 : boolean;
  signal addr_of_3426_final_reg_ack_1 : boolean;
  signal type_cast_3095_inst_req_0 : boolean;
  signal type_cast_3095_inst_ack_0 : boolean;
  signal type_cast_3095_inst_req_1 : boolean;
  signal type_cast_3095_inst_ack_1 : boolean;
  signal type_cast_3164_inst_req_0 : boolean;
  signal type_cast_3164_inst_ack_0 : boolean;
  signal type_cast_3164_inst_req_1 : boolean;
  signal type_cast_3164_inst_ack_1 : boolean;
  signal if_stmt_3173_branch_req_0 : boolean;
  signal type_cast_3605_inst_ack_0 : boolean;
  signal if_stmt_3173_branch_ack_1 : boolean;
  signal if_stmt_3173_branch_ack_0 : boolean;
  signal type_cast_3483_inst_ack_1 : boolean;
  signal type_cast_3483_inst_req_1 : boolean;
  signal LOAD_row_high_3181_load_0_req_0 : boolean;
  signal LOAD_row_high_3181_load_0_ack_0 : boolean;
  signal type_cast_3437_inst_ack_1 : boolean;
  signal LOAD_row_high_3181_load_0_req_1 : boolean;
  signal LOAD_row_high_3181_load_0_ack_1 : boolean;
  signal type_cast_3605_inst_req_0 : boolean;
  signal type_cast_3476_inst_ack_1 : boolean;
  signal type_cast_3476_inst_req_1 : boolean;
  signal if_stmt_3551_branch_ack_0 : boolean;
  signal type_cast_3185_inst_req_0 : boolean;
  signal type_cast_3185_inst_ack_0 : boolean;
  signal addr_of_3426_final_reg_req_1 : boolean;
  signal type_cast_3185_inst_req_1 : boolean;
  signal type_cast_3185_inst_ack_1 : boolean;
  signal type_cast_4095_inst_req_1 : boolean;
  signal LOAD_row_high_3523_load_0_ack_1 : boolean;
  signal type_cast_3527_inst_ack_0 : boolean;
  signal ptr_deref_3429_store_0_ack_1 : boolean;
  signal if_stmt_3551_branch_ack_1 : boolean;
  signal if_stmt_3211_branch_req_0 : boolean;
  signal type_cast_3476_inst_ack_0 : boolean;
  signal ptr_deref_4011_store_0_ack_0 : boolean;
  signal if_stmt_3211_branch_ack_1 : boolean;
  signal if_stmt_3211_branch_ack_0 : boolean;
  signal type_cast_3483_inst_ack_0 : boolean;
  signal type_cast_3483_inst_req_0 : boolean;
  signal type_cast_3476_inst_req_0 : boolean;
  signal type_cast_3221_inst_req_0 : boolean;
  signal type_cast_3221_inst_ack_0 : boolean;
  signal type_cast_3520_inst_ack_1 : boolean;
  signal type_cast_3221_inst_req_1 : boolean;
  signal type_cast_3221_inst_ack_1 : boolean;
  signal type_cast_3520_inst_req_1 : boolean;
  signal if_stmt_3230_branch_req_0 : boolean;
  signal if_stmt_3230_branch_ack_1 : boolean;
  signal addr_of_3426_final_reg_ack_0 : boolean;
  signal if_stmt_3230_branch_ack_0 : boolean;
  signal type_cast_3527_inst_req_0 : boolean;
  signal type_cast_3437_inst_req_1 : boolean;
  signal LOAD_col_high_3238_load_0_req_0 : boolean;
  signal LOAD_col_high_3238_load_0_ack_0 : boolean;
  signal LOAD_col_high_3238_load_0_req_1 : boolean;
  signal LOAD_col_high_3238_load_0_ack_1 : boolean;
  signal if_stmt_3452_branch_ack_0 : boolean;
  signal type_cast_3520_inst_ack_0 : boolean;
  signal type_cast_3242_inst_req_0 : boolean;
  signal type_cast_3520_inst_req_0 : boolean;
  signal type_cast_3242_inst_ack_0 : boolean;
  signal addr_of_3426_final_reg_req_0 : boolean;
  signal if_stmt_3551_branch_req_0 : boolean;
  signal type_cast_3242_inst_req_1 : boolean;
  signal type_cast_3242_inst_ack_1 : boolean;
  signal ptr_deref_3429_store_0_req_1 : boolean;
  signal LOAD_row_high_3523_load_0_req_1 : boolean;
  signal if_stmt_3262_branch_req_0 : boolean;
  signal if_stmt_3452_branch_ack_1 : boolean;
  signal if_stmt_3262_branch_ack_1 : boolean;
  signal if_stmt_3262_branch_ack_0 : boolean;
  signal type_cast_3272_inst_req_0 : boolean;
  signal type_cast_3272_inst_ack_0 : boolean;
  signal type_cast_3272_inst_req_1 : boolean;
  signal type_cast_3272_inst_ack_1 : boolean;
  signal type_cast_4095_inst_ack_1 : boolean;
  signal type_cast_4065_inst_ack_0 : boolean;
  signal type_cast_3277_inst_req_0 : boolean;
  signal type_cast_3277_inst_ack_0 : boolean;
  signal type_cast_3277_inst_req_1 : boolean;
  signal type_cast_3277_inst_ack_1 : boolean;
  signal type_cast_3311_inst_req_0 : boolean;
  signal type_cast_3311_inst_ack_0 : boolean;
  signal type_cast_3311_inst_req_1 : boolean;
  signal type_cast_3311_inst_ack_1 : boolean;
  signal type_cast_4019_inst_req_1 : boolean;
  signal array_obj_ref_3317_index_offset_req_0 : boolean;
  signal array_obj_ref_3317_index_offset_ack_0 : boolean;
  signal array_obj_ref_3317_index_offset_req_1 : boolean;
  signal if_stmt_4126_branch_req_0 : boolean;
  signal array_obj_ref_3317_index_offset_ack_1 : boolean;
  signal type_cast_4019_inst_ack_1 : boolean;
  signal type_cast_4065_inst_req_1 : boolean;
  signal addr_of_3318_final_reg_req_0 : boolean;
  signal addr_of_3318_final_reg_ack_0 : boolean;
  signal addr_of_3318_final_reg_req_1 : boolean;
  signal addr_of_3318_final_reg_ack_1 : boolean;
  signal type_cast_4065_inst_ack_1 : boolean;
  signal ptr_deref_3321_store_0_req_0 : boolean;
  signal ptr_deref_3321_store_0_ack_0 : boolean;
  signal ptr_deref_3321_store_0_req_1 : boolean;
  signal ptr_deref_3321_store_0_ack_1 : boolean;
  signal LOAD_pad_4181_load_0_ack_1 : boolean;
  signal type_cast_3330_inst_req_0 : boolean;
  signal type_cast_3330_inst_ack_0 : boolean;
  signal type_cast_3330_inst_req_1 : boolean;
  signal type_cast_3330_inst_ack_1 : boolean;
  signal type_cast_3394_inst_req_0 : boolean;
  signal type_cast_3394_inst_ack_0 : boolean;
  signal type_cast_3394_inst_req_1 : boolean;
  signal if_stmt_4126_branch_ack_1 : boolean;
  signal type_cast_3394_inst_ack_1 : boolean;
  signal if_stmt_4034_branch_req_0 : boolean;
  signal array_obj_ref_3400_index_offset_req_0 : boolean;
  signal array_obj_ref_3400_index_offset_ack_0 : boolean;
  signal array_obj_ref_3400_index_offset_req_1 : boolean;
  signal array_obj_ref_3400_index_offset_ack_1 : boolean;
  signal addr_of_3401_final_reg_req_0 : boolean;
  signal addr_of_3401_final_reg_ack_0 : boolean;
  signal addr_of_3401_final_reg_req_1 : boolean;
  signal addr_of_3401_final_reg_ack_1 : boolean;
  signal ptr_deref_3405_load_0_req_0 : boolean;
  signal ptr_deref_3405_load_0_ack_0 : boolean;
  signal ptr_deref_3405_load_0_req_1 : boolean;
  signal ptr_deref_3405_load_0_ack_1 : boolean;
  signal type_cast_3419_inst_req_0 : boolean;
  signal type_cast_3419_inst_ack_0 : boolean;
  signal type_cast_3419_inst_req_1 : boolean;
  signal type_cast_3419_inst_ack_1 : boolean;
  signal array_obj_ref_3425_index_offset_req_0 : boolean;
  signal array_obj_ref_3425_index_offset_ack_0 : boolean;
  signal array_obj_ref_3425_index_offset_req_1 : boolean;
  signal array_obj_ref_3425_index_offset_ack_1 : boolean;
  signal LOAD_pad_3614_load_0_req_0 : boolean;
  signal LOAD_pad_3614_load_0_ack_0 : boolean;
  signal LOAD_pad_3614_load_0_req_1 : boolean;
  signal LOAD_pad_3614_load_0_ack_1 : boolean;
  signal LOAD_depth_high_3617_load_0_req_0 : boolean;
  signal LOAD_depth_high_3617_load_0_ack_0 : boolean;
  signal LOAD_depth_high_3617_load_0_req_1 : boolean;
  signal LOAD_depth_high_3617_load_0_ack_1 : boolean;
  signal ptr_deref_3629_load_0_req_0 : boolean;
  signal ptr_deref_3629_load_0_ack_0 : boolean;
  signal ptr_deref_3629_load_0_req_1 : boolean;
  signal ptr_deref_3629_load_0_ack_1 : boolean;
  signal ptr_deref_3641_load_0_req_0 : boolean;
  signal ptr_deref_3641_load_0_ack_0 : boolean;
  signal ptr_deref_3641_load_0_req_1 : boolean;
  signal ptr_deref_3641_load_0_ack_1 : boolean;
  signal type_cast_3645_inst_req_0 : boolean;
  signal type_cast_3645_inst_ack_0 : boolean;
  signal type_cast_3645_inst_req_1 : boolean;
  signal type_cast_3645_inst_ack_1 : boolean;
  signal type_cast_3684_inst_req_0 : boolean;
  signal type_cast_3684_inst_ack_0 : boolean;
  signal type_cast_3684_inst_req_1 : boolean;
  signal type_cast_3684_inst_ack_1 : boolean;
  signal type_cast_3752_inst_req_0 : boolean;
  signal type_cast_3752_inst_ack_0 : boolean;
  signal type_cast_3752_inst_req_1 : boolean;
  signal type_cast_3752_inst_ack_1 : boolean;
  signal if_stmt_3761_branch_req_0 : boolean;
  signal if_stmt_3761_branch_ack_1 : boolean;
  signal if_stmt_3761_branch_ack_0 : boolean;
  signal LOAD_row_high_3769_load_0_req_0 : boolean;
  signal LOAD_row_high_3769_load_0_ack_0 : boolean;
  signal ptr_deref_4011_store_0_req_0 : boolean;
  signal LOAD_row_high_3769_load_0_req_1 : boolean;
  signal LOAD_row_high_3769_load_0_ack_1 : boolean;
  signal type_cast_4019_inst_ack_0 : boolean;
  signal type_cast_4065_inst_req_0 : boolean;
  signal type_cast_3773_inst_req_0 : boolean;
  signal type_cast_4102_inst_ack_1 : boolean;
  signal type_cast_3773_inst_ack_0 : boolean;
  signal type_cast_3773_inst_req_1 : boolean;
  signal type_cast_4102_inst_req_1 : boolean;
  signal type_cast_3773_inst_ack_1 : boolean;
  signal if_stmt_3799_branch_req_0 : boolean;
  signal type_cast_4095_inst_ack_0 : boolean;
  signal if_stmt_3799_branch_ack_1 : boolean;
  signal type_cast_4095_inst_req_0 : boolean;
  signal if_stmt_3799_branch_ack_0 : boolean;
  signal type_cast_3809_inst_req_0 : boolean;
  signal type_cast_3809_inst_ack_0 : boolean;
  signal type_cast_4102_inst_ack_0 : boolean;
  signal type_cast_3809_inst_req_1 : boolean;
  signal type_cast_3809_inst_ack_1 : boolean;
  signal type_cast_4019_inst_req_0 : boolean;
  signal LOAD_depth_high_4184_load_0_ack_1 : boolean;
  signal if_stmt_3818_branch_req_0 : boolean;
  signal if_stmt_3818_branch_ack_1 : boolean;
  signal if_stmt_3818_branch_ack_0 : boolean;
  signal type_cast_4102_inst_req_0 : boolean;
  signal LOAD_pad_4181_load_0_req_1 : boolean;
  signal LOAD_depth_high_4184_load_0_req_1 : boolean;
  signal LOAD_col_high_3826_load_0_req_0 : boolean;
  signal LOAD_col_high_3826_load_0_ack_0 : boolean;
  signal if_stmt_4034_branch_ack_0 : boolean;
  signal LOAD_col_high_3826_load_0_req_1 : boolean;
  signal LOAD_col_high_3826_load_0_ack_1 : boolean;
  signal type_cast_4079_inst_ack_1 : boolean;
  signal LOAD_col_high_4061_load_0_ack_1 : boolean;
  signal type_cast_3830_inst_req_0 : boolean;
  signal type_cast_3830_inst_ack_0 : boolean;
  signal type_cast_4079_inst_req_1 : boolean;
  signal type_cast_3830_inst_req_1 : boolean;
  signal type_cast_3830_inst_ack_1 : boolean;
  signal ptr_deref_4196_load_0_ack_0 : boolean;
  signal LOAD_col_high_4061_load_0_req_1 : boolean;
  signal if_stmt_3844_branch_req_0 : boolean;
  signal if_stmt_3844_branch_ack_1 : boolean;
  signal type_cast_4079_inst_ack_0 : boolean;
  signal if_stmt_3844_branch_ack_0 : boolean;
  signal LOAD_pad_4181_load_0_ack_0 : boolean;
  signal type_cast_4079_inst_req_0 : boolean;
  signal type_cast_3854_inst_req_0 : boolean;
  signal type_cast_3854_inst_ack_0 : boolean;
  signal LOAD_depth_high_4184_load_0_ack_0 : boolean;
  signal LOAD_depth_high_4184_load_0_req_0 : boolean;
  signal type_cast_3854_inst_req_1 : boolean;
  signal type_cast_3854_inst_ack_1 : boolean;
  signal ptr_deref_4196_load_0_req_0 : boolean;
  signal addr_of_4008_final_reg_ack_1 : boolean;
  signal type_cast_3859_inst_req_0 : boolean;
  signal type_cast_3859_inst_ack_0 : boolean;
  signal type_cast_3859_inst_req_1 : boolean;
  signal type_cast_3859_inst_ack_1 : boolean;
  signal type_cast_3893_inst_req_0 : boolean;
  signal type_cast_3893_inst_ack_0 : boolean;
  signal type_cast_3893_inst_req_1 : boolean;
  signal type_cast_3893_inst_ack_1 : boolean;
  signal type_cast_4166_inst_ack_1 : boolean;
  signal type_cast_4166_inst_req_1 : boolean;
  signal type_cast_4166_inst_ack_0 : boolean;
  signal addr_of_4008_final_reg_req_1 : boolean;
  signal LOAD_col_high_4061_load_0_ack_0 : boolean;
  signal array_obj_ref_3899_index_offset_req_0 : boolean;
  signal LOAD_row_high_4098_load_0_ack_1 : boolean;
  signal array_obj_ref_3899_index_offset_ack_0 : boolean;
  signal array_obj_ref_3899_index_offset_req_1 : boolean;
  signal LOAD_row_high_4098_load_0_req_1 : boolean;
  signal array_obj_ref_3899_index_offset_ack_1 : boolean;
  signal LOAD_col_high_4061_load_0_req_0 : boolean;
  signal addr_of_3900_final_reg_req_0 : boolean;
  signal addr_of_3900_final_reg_ack_0 : boolean;
  signal addr_of_3900_final_reg_req_1 : boolean;
  signal addr_of_3900_final_reg_ack_1 : boolean;
  signal type_cast_4166_inst_req_0 : boolean;
  signal LOAD_row_high_4098_load_0_ack_0 : boolean;
  signal LOAD_row_high_4098_load_0_req_0 : boolean;
  signal if_stmt_4034_branch_ack_1 : boolean;
  signal ptr_deref_3903_store_0_req_0 : boolean;
  signal ptr_deref_3903_store_0_ack_0 : boolean;
  signal addr_of_4008_final_reg_ack_0 : boolean;
  signal ptr_deref_3903_store_0_req_1 : boolean;
  signal ptr_deref_3903_store_0_ack_1 : boolean;
  signal addr_of_4008_final_reg_req_0 : boolean;
  signal type_cast_4620_inst_req_0 : boolean;
  signal type_cast_3912_inst_req_0 : boolean;
  signal type_cast_3912_inst_ack_0 : boolean;
  signal type_cast_3912_inst_req_1 : boolean;
  signal type_cast_3912_inst_ack_1 : boolean;
  signal ptr_deref_4011_store_0_ack_1 : boolean;
  signal if_stmt_4126_branch_ack_0 : boolean;
  signal LOAD_pad_4181_load_0_req_0 : boolean;
  signal type_cast_3976_inst_req_0 : boolean;
  signal type_cast_3976_inst_ack_0 : boolean;
  signal type_cast_3976_inst_req_1 : boolean;
  signal type_cast_3976_inst_ack_1 : boolean;
  signal ptr_deref_4011_store_0_req_1 : boolean;
  signal type_cast_4058_inst_ack_1 : boolean;
  signal type_cast_4058_inst_req_1 : boolean;
  signal type_cast_4058_inst_ack_0 : boolean;
  signal type_cast_4058_inst_req_0 : boolean;
  signal array_obj_ref_3982_index_offset_req_0 : boolean;
  signal array_obj_ref_3982_index_offset_ack_0 : boolean;
  signal array_obj_ref_3982_index_offset_req_1 : boolean;
  signal array_obj_ref_3982_index_offset_ack_1 : boolean;
  signal addr_of_3983_final_reg_req_0 : boolean;
  signal addr_of_3983_final_reg_ack_0 : boolean;
  signal addr_of_3983_final_reg_req_1 : boolean;
  signal type_cast_4664_inst_req_1 : boolean;
  signal addr_of_3983_final_reg_ack_1 : boolean;
  signal type_cast_4664_inst_ack_1 : boolean;
  signal ptr_deref_3987_load_0_req_0 : boolean;
  signal ptr_deref_3987_load_0_ack_0 : boolean;
  signal LOAD_col_high_4623_load_0_ack_0 : boolean;
  signal ptr_deref_3987_load_0_req_1 : boolean;
  signal ptr_deref_3987_load_0_ack_1 : boolean;
  signal type_cast_4001_inst_req_0 : boolean;
  signal type_cast_4001_inst_ack_0 : boolean;
  signal type_cast_4001_inst_req_1 : boolean;
  signal type_cast_4001_inst_ack_1 : boolean;
  signal array_obj_ref_4007_index_offset_req_0 : boolean;
  signal array_obj_ref_4007_index_offset_ack_0 : boolean;
  signal array_obj_ref_4007_index_offset_req_1 : boolean;
  signal array_obj_ref_4007_index_offset_ack_1 : boolean;
  signal ptr_deref_4196_load_0_req_1 : boolean;
  signal ptr_deref_4196_load_0_ack_1 : boolean;
  signal ptr_deref_4208_load_0_req_0 : boolean;
  signal ptr_deref_4208_load_0_ack_0 : boolean;
  signal ptr_deref_4208_load_0_req_1 : boolean;
  signal ptr_deref_4208_load_0_ack_1 : boolean;
  signal type_cast_4212_inst_req_0 : boolean;
  signal type_cast_4212_inst_ack_0 : boolean;
  signal type_cast_4212_inst_req_1 : boolean;
  signal type_cast_4212_inst_ack_1 : boolean;
  signal type_cast_4251_inst_req_0 : boolean;
  signal type_cast_4251_inst_ack_0 : boolean;
  signal type_cast_4251_inst_req_1 : boolean;
  signal type_cast_4251_inst_ack_1 : boolean;
  signal type_cast_4320_inst_req_0 : boolean;
  signal type_cast_4320_inst_ack_0 : boolean;
  signal type_cast_4320_inst_req_1 : boolean;
  signal type_cast_4320_inst_ack_1 : boolean;
  signal if_stmt_4329_branch_req_0 : boolean;
  signal if_stmt_4329_branch_ack_1 : boolean;
  signal if_stmt_4329_branch_ack_0 : boolean;
  signal LOAD_row_high_4337_load_0_req_0 : boolean;
  signal LOAD_row_high_4337_load_0_ack_0 : boolean;
  signal LOAD_row_high_4337_load_0_req_1 : boolean;
  signal LOAD_row_high_4337_load_0_ack_1 : boolean;
  signal type_cast_4341_inst_req_0 : boolean;
  signal type_cast_4341_inst_ack_0 : boolean;
  signal type_cast_4341_inst_req_1 : boolean;
  signal type_cast_4341_inst_ack_1 : boolean;
  signal type_cast_4822_inst_ack_0 : boolean;
  signal type_cast_4783_inst_ack_1 : boolean;
  signal type_cast_4664_inst_ack_0 : boolean;
  signal if_stmt_4355_branch_req_0 : boolean;
  signal type_cast_4822_inst_req_0 : boolean;
  signal if_stmt_4355_branch_ack_1 : boolean;
  signal if_stmt_4355_branch_ack_0 : boolean;
  signal type_cast_4365_inst_req_0 : boolean;
  signal type_cast_4365_inst_ack_0 : boolean;
  signal type_cast_4737_inst_ack_1 : boolean;
  signal type_cast_4365_inst_req_1 : boolean;
  signal type_cast_4365_inst_ack_1 : boolean;
  signal type_cast_4737_inst_req_1 : boolean;
  signal if_stmt_4596_branch_ack_0 : boolean;
  signal if_stmt_4374_branch_req_0 : boolean;
  signal if_stmt_4596_branch_ack_1 : boolean;
  signal if_stmt_4374_branch_ack_1 : boolean;
  signal if_stmt_4374_branch_ack_0 : boolean;
  signal type_cast_4783_inst_req_1 : boolean;
  signal type_cast_4664_inst_req_0 : boolean;
  signal LOAD_col_high_4623_load_0_req_0 : boolean;
  signal LOAD_col_high_4382_load_0_req_0 : boolean;
  signal LOAD_col_high_4382_load_0_ack_0 : boolean;
  signal LOAD_col_high_4382_load_0_req_1 : boolean;
  signal LOAD_col_high_4382_load_0_ack_1 : boolean;
  signal LOAD_row_high_4667_load_0_ack_1 : boolean;
  signal type_cast_4890_inst_req_1 : boolean;
  signal ptr_deref_4779_load_0_ack_0 : boolean;
  signal type_cast_4737_inst_ack_0 : boolean;
  signal type_cast_4386_inst_req_0 : boolean;
  signal type_cast_4737_inst_req_0 : boolean;
  signal type_cast_4386_inst_ack_0 : boolean;
  signal LOAD_row_high_4667_load_0_req_1 : boolean;
  signal type_cast_4386_inst_req_1 : boolean;
  signal type_cast_4386_inst_ack_1 : boolean;
  signal type_cast_4890_inst_ack_0 : boolean;
  signal type_cast_4647_inst_ack_1 : boolean;
  signal if_stmt_4406_branch_req_0 : boolean;
  signal ptr_deref_4779_load_0_req_0 : boolean;
  signal type_cast_4647_inst_req_1 : boolean;
  signal if_stmt_4596_branch_req_0 : boolean;
  signal if_stmt_4406_branch_ack_1 : boolean;
  signal if_stmt_4406_branch_ack_0 : boolean;
  signal type_cast_4416_inst_req_0 : boolean;
  signal type_cast_4416_inst_ack_0 : boolean;
  signal type_cast_4416_inst_req_1 : boolean;
  signal type_cast_4416_inst_ack_1 : boolean;
  signal type_cast_4581_inst_ack_1 : boolean;
  signal type_cast_4421_inst_req_0 : boolean;
  signal type_cast_4421_inst_ack_0 : boolean;
  signal type_cast_4421_inst_req_1 : boolean;
  signal type_cast_4421_inst_ack_1 : boolean;
  signal type_cast_4581_inst_req_1 : boolean;
  signal type_cast_4890_inst_ack_1 : boolean;
  signal type_cast_4783_inst_ack_0 : boolean;
  signal type_cast_4455_inst_req_0 : boolean;
  signal type_cast_4727_inst_ack_1 : boolean;
  signal type_cast_4455_inst_ack_0 : boolean;
  signal type_cast_4455_inst_req_1 : boolean;
  signal type_cast_4727_inst_req_1 : boolean;
  signal type_cast_4455_inst_ack_1 : boolean;
  signal type_cast_4783_inst_req_0 : boolean;
  signal type_cast_4890_inst_req_0 : boolean;
  signal type_cast_4647_inst_ack_0 : boolean;
  signal type_cast_4647_inst_req_0 : boolean;
  signal LOAD_row_high_4667_load_0_ack_0 : boolean;
  signal array_obj_ref_4461_index_offset_req_0 : boolean;
  signal array_obj_ref_4461_index_offset_ack_0 : boolean;
  signal array_obj_ref_4461_index_offset_req_1 : boolean;
  signal array_obj_ref_4461_index_offset_ack_1 : boolean;
  signal type_cast_4727_inst_ack_0 : boolean;
  signal type_cast_4620_inst_ack_1 : boolean;
  signal type_cast_4727_inst_req_0 : boolean;
  signal addr_of_4462_final_reg_req_0 : boolean;
  signal addr_of_4462_final_reg_ack_0 : boolean;
  signal LOAD_row_high_4667_load_0_req_0 : boolean;
  signal addr_of_4462_final_reg_req_1 : boolean;
  signal addr_of_4462_final_reg_ack_1 : boolean;
  signal type_cast_4822_inst_req_1 : boolean;
  signal LOAD_depth_high_4755_load_0_ack_1 : boolean;
  signal LOAD_depth_high_4755_load_0_req_1 : boolean;
  signal ptr_deref_4465_store_0_req_0 : boolean;
  signal type_cast_4627_inst_ack_1 : boolean;
  signal ptr_deref_4465_store_0_ack_0 : boolean;
  signal type_cast_4581_inst_ack_0 : boolean;
  signal ptr_deref_4465_store_0_req_1 : boolean;
  signal ptr_deref_4465_store_0_ack_1 : boolean;
  signal type_cast_4581_inst_req_0 : boolean;
  signal type_cast_4627_inst_req_1 : boolean;
  signal ptr_deref_4767_load_0_ack_1 : boolean;
  signal type_cast_4474_inst_req_0 : boolean;
  signal type_cast_4474_inst_ack_0 : boolean;
  signal ptr_deref_4767_load_0_req_1 : boolean;
  signal type_cast_4474_inst_req_1 : boolean;
  signal if_stmt_4683_branch_ack_0 : boolean;
  signal type_cast_4474_inst_ack_1 : boolean;
  signal ptr_deref_4573_store_0_ack_1 : boolean;
  signal type_cast_4538_inst_req_0 : boolean;
  signal type_cast_4538_inst_ack_0 : boolean;
  signal type_cast_4538_inst_req_1 : boolean;
  signal type_cast_4538_inst_ack_1 : boolean;
  signal LOAD_depth_high_4755_load_0_ack_0 : boolean;
  signal LOAD_depth_high_4755_load_0_req_0 : boolean;
  signal type_cast_4627_inst_ack_0 : boolean;
  signal ptr_deref_4573_store_0_req_1 : boolean;
  signal type_cast_4627_inst_req_0 : boolean;
  signal array_obj_ref_4544_index_offset_req_0 : boolean;
  signal if_stmt_4683_branch_ack_1 : boolean;
  signal array_obj_ref_4544_index_offset_ack_0 : boolean;
  signal type_cast_4620_inst_req_1 : boolean;
  signal array_obj_ref_4544_index_offset_req_1 : boolean;
  signal array_obj_ref_4544_index_offset_ack_1 : boolean;
  signal if_stmt_4683_branch_req_0 : boolean;
  signal addr_of_4545_final_reg_req_0 : boolean;
  signal addr_of_4545_final_reg_ack_0 : boolean;
  signal addr_of_4545_final_reg_req_1 : boolean;
  signal addr_of_4545_final_reg_ack_1 : boolean;
  signal type_cast_4671_inst_ack_1 : boolean;
  signal ptr_deref_4549_load_0_req_0 : boolean;
  signal ptr_deref_4549_load_0_ack_0 : boolean;
  signal ptr_deref_4549_load_0_req_1 : boolean;
  signal ptr_deref_4549_load_0_ack_1 : boolean;
  signal ptr_deref_4767_load_0_ack_0 : boolean;
  signal ptr_deref_4779_load_0_ack_1 : boolean;
  signal ptr_deref_4779_load_0_req_1 : boolean;
  signal LOAD_col_high_4623_load_0_ack_1 : boolean;
  signal ptr_deref_4767_load_0_req_0 : boolean;
  signal LOAD_col_high_4623_load_0_req_1 : boolean;
  signal type_cast_4563_inst_req_0 : boolean;
  signal type_cast_4671_inst_req_1 : boolean;
  signal type_cast_4563_inst_ack_0 : boolean;
  signal type_cast_4563_inst_req_1 : boolean;
  signal type_cast_4563_inst_ack_1 : boolean;
  signal LOAD_pad_4752_load_0_ack_1 : boolean;
  signal LOAD_pad_4752_load_0_req_1 : boolean;
  signal array_obj_ref_4569_index_offset_req_0 : boolean;
  signal array_obj_ref_4569_index_offset_ack_0 : boolean;
  signal type_cast_4620_inst_ack_0 : boolean;
  signal array_obj_ref_4569_index_offset_req_1 : boolean;
  signal type_cast_4671_inst_ack_0 : boolean;
  signal array_obj_ref_4569_index_offset_ack_1 : boolean;
  signal type_cast_4822_inst_ack_1 : boolean;
  signal type_cast_4671_inst_req_0 : boolean;
  signal addr_of_4570_final_reg_req_0 : boolean;
  signal addr_of_4570_final_reg_ack_0 : boolean;
  signal addr_of_4570_final_reg_req_1 : boolean;
  signal addr_of_4570_final_reg_ack_1 : boolean;
  signal LOAD_pad_4752_load_0_ack_0 : boolean;
  signal LOAD_pad_4752_load_0_req_0 : boolean;
  signal ptr_deref_4573_store_0_req_0 : boolean;
  signal ptr_deref_4573_store_0_ack_0 : boolean;
  signal if_stmt_4899_branch_req_0 : boolean;
  signal if_stmt_4899_branch_ack_1 : boolean;
  signal if_stmt_4899_branch_ack_0 : boolean;
  signal LOAD_row_high_4907_load_0_req_0 : boolean;
  signal LOAD_row_high_4907_load_0_ack_0 : boolean;
  signal LOAD_row_high_4907_load_0_req_1 : boolean;
  signal LOAD_row_high_4907_load_0_ack_1 : boolean;
  signal type_cast_4911_inst_req_0 : boolean;
  signal type_cast_4911_inst_ack_0 : boolean;
  signal type_cast_4911_inst_req_1 : boolean;
  signal type_cast_4911_inst_ack_1 : boolean;
  signal if_stmt_4925_branch_req_0 : boolean;
  signal if_stmt_4925_branch_ack_1 : boolean;
  signal if_stmt_4925_branch_ack_0 : boolean;
  signal type_cast_4935_inst_req_0 : boolean;
  signal type_cast_4935_inst_ack_0 : boolean;
  signal type_cast_4935_inst_req_1 : boolean;
  signal type_cast_4935_inst_ack_1 : boolean;
  signal if_stmt_4944_branch_req_0 : boolean;
  signal if_stmt_4944_branch_ack_1 : boolean;
  signal if_stmt_4944_branch_ack_0 : boolean;
  signal type_cast_1312_inst_ack_1 : boolean;
  signal phi_stmt_899_req_1 : boolean;
  signal type_cast_1318_inst_req_1 : boolean;
  signal type_cast_905_inst_ack_1 : boolean;
  signal LOAD_col_high_4952_load_0_req_0 : boolean;
  signal type_cast_905_inst_req_1 : boolean;
  signal LOAD_col_high_4952_load_0_ack_0 : boolean;
  signal LOAD_col_high_4952_load_0_req_1 : boolean;
  signal LOAD_col_high_4952_load_0_ack_1 : boolean;
  signal type_cast_905_inst_ack_0 : boolean;
  signal type_cast_1325_inst_req_0 : boolean;
  signal type_cast_905_inst_req_0 : boolean;
  signal type_cast_4956_inst_req_0 : boolean;
  signal type_cast_4956_inst_ack_0 : boolean;
  signal phi_stmt_906_req_1 : boolean;
  signal type_cast_4956_inst_req_1 : boolean;
  signal type_cast_4956_inst_ack_1 : boolean;
  signal type_cast_1312_inst_req_1 : boolean;
  signal type_cast_912_inst_ack_1 : boolean;
  signal if_stmt_4970_branch_req_0 : boolean;
  signal type_cast_912_inst_req_1 : boolean;
  signal LOAD_row_high_5224_load_0_ack_1 : boolean;
  signal if_stmt_4970_branch_ack_1 : boolean;
  signal LOAD_row_high_5224_load_0_req_1 : boolean;
  signal if_stmt_4970_branch_ack_0 : boolean;
  signal type_cast_1318_inst_req_0 : boolean;
  signal if_stmt_5240_branch_req_0 : boolean;
  signal type_cast_4980_inst_req_0 : boolean;
  signal type_cast_4980_inst_ack_0 : boolean;
  signal type_cast_4980_inst_req_1 : boolean;
  signal type_cast_4980_inst_ack_1 : boolean;
  signal phi_stmt_1307_req_0 : boolean;
  signal type_cast_4985_inst_req_0 : boolean;
  signal type_cast_4985_inst_ack_0 : boolean;
  signal type_cast_1310_inst_ack_1 : boolean;
  signal type_cast_4985_inst_req_1 : boolean;
  signal type_cast_4985_inst_ack_1 : boolean;
  signal type_cast_1312_inst_ack_0 : boolean;
  signal type_cast_1312_inst_req_0 : boolean;
  signal type_cast_1310_inst_req_1 : boolean;
  signal type_cast_5019_inst_req_0 : boolean;
  signal type_cast_5019_inst_ack_0 : boolean;
  signal type_cast_1310_inst_ack_0 : boolean;
  signal type_cast_5019_inst_req_1 : boolean;
  signal type_cast_5019_inst_ack_1 : boolean;
  signal type_cast_1310_inst_req_0 : boolean;
  signal type_cast_912_inst_ack_0 : boolean;
  signal type_cast_912_inst_req_0 : boolean;
  signal array_obj_ref_5025_index_offset_req_0 : boolean;
  signal array_obj_ref_5025_index_offset_ack_0 : boolean;
  signal array_obj_ref_5025_index_offset_req_1 : boolean;
  signal array_obj_ref_5025_index_offset_ack_1 : boolean;
  signal type_cast_5228_inst_ack_0 : boolean;
  signal phi_stmt_1313_req_0 : boolean;
  signal addr_of_5026_final_reg_req_0 : boolean;
  signal addr_of_5026_final_reg_ack_0 : boolean;
  signal addr_of_5026_final_reg_req_1 : boolean;
  signal addr_of_5026_final_reg_ack_1 : boolean;
  signal phi_stmt_913_req_0 : boolean;
  signal ptr_deref_5029_store_0_req_0 : boolean;
  signal ptr_deref_5029_store_0_ack_0 : boolean;
  signal LOAD_row_high_5224_load_0_ack_0 : boolean;
  signal ptr_deref_5029_store_0_req_1 : boolean;
  signal ptr_deref_5029_store_0_ack_1 : boolean;
  signal LOAD_row_high_5224_load_0_req_0 : boolean;
  signal type_cast_1316_inst_ack_1 : boolean;
  signal type_cast_1316_inst_req_1 : boolean;
  signal type_cast_5038_inst_req_0 : boolean;
  signal type_cast_5038_inst_ack_0 : boolean;
  signal type_cast_5038_inst_req_1 : boolean;
  signal type_cast_5038_inst_ack_1 : boolean;
  signal type_cast_5102_inst_req_0 : boolean;
  signal type_cast_5102_inst_ack_0 : boolean;
  signal type_cast_5102_inst_req_1 : boolean;
  signal type_cast_5102_inst_ack_1 : boolean;
  signal phi_stmt_906_req_0 : boolean;
  signal array_obj_ref_5108_index_offset_req_0 : boolean;
  signal array_obj_ref_5108_index_offset_ack_0 : boolean;
  signal type_cast_5228_inst_req_0 : boolean;
  signal array_obj_ref_5108_index_offset_req_1 : boolean;
  signal array_obj_ref_5108_index_offset_ack_1 : boolean;
  signal type_cast_1316_inst_ack_0 : boolean;
  signal phi_stmt_913_ack_0 : boolean;
  signal addr_of_5109_final_reg_req_0 : boolean;
  signal phi_stmt_906_ack_0 : boolean;
  signal addr_of_5109_final_reg_ack_0 : boolean;
  signal phi_stmt_1319_req_0 : boolean;
  signal addr_of_5109_final_reg_req_1 : boolean;
  signal phi_stmt_899_ack_0 : boolean;
  signal addr_of_5109_final_reg_ack_1 : boolean;
  signal phi_stmt_1319_req_1 : boolean;
  signal type_cast_1325_inst_ack_1 : boolean;
  signal phi_stmt_899_req_0 : boolean;
  signal phi_stmt_913_req_1 : boolean;
  signal ptr_deref_5113_load_0_req_0 : boolean;
  signal ptr_deref_5113_load_0_ack_0 : boolean;
  signal type_cast_5228_inst_ack_1 : boolean;
  signal ptr_deref_5113_load_0_req_1 : boolean;
  signal ptr_deref_5113_load_0_ack_1 : boolean;
  signal type_cast_1325_inst_req_1 : boolean;
  signal type_cast_1318_inst_ack_0 : boolean;
  signal type_cast_5127_inst_req_0 : boolean;
  signal type_cast_919_inst_ack_1 : boolean;
  signal type_cast_5127_inst_ack_0 : boolean;
  signal type_cast_5127_inst_req_1 : boolean;
  signal type_cast_919_inst_req_1 : boolean;
  signal type_cast_5127_inst_ack_1 : boolean;
  signal type_cast_1325_inst_ack_0 : boolean;
  signal call_stmt_5270_call_ack_1 : boolean;
  signal call_stmt_5270_call_req_1 : boolean;
  signal array_obj_ref_5133_index_offset_req_0 : boolean;
  signal array_obj_ref_5133_index_offset_ack_0 : boolean;
  signal array_obj_ref_5133_index_offset_req_1 : boolean;
  signal array_obj_ref_5133_index_offset_ack_1 : boolean;
  signal type_cast_1316_inst_req_0 : boolean;
  signal call_stmt_5270_call_ack_0 : boolean;
  signal type_cast_919_inst_ack_0 : boolean;
  signal type_cast_919_inst_req_0 : boolean;
  signal addr_of_5134_final_reg_req_0 : boolean;
  signal addr_of_5134_final_reg_ack_0 : boolean;
  signal phi_stmt_1313_req_1 : boolean;
  signal addr_of_5134_final_reg_req_1 : boolean;
  signal addr_of_5134_final_reg_ack_1 : boolean;
  signal call_stmt_5270_call_req_0 : boolean;
  signal if_stmt_5240_branch_ack_0 : boolean;
  signal type_cast_5221_inst_ack_1 : boolean;
  signal type_cast_5228_inst_req_1 : boolean;
  signal type_cast_1318_inst_ack_1 : boolean;
  signal if_stmt_5240_branch_ack_1 : boolean;
  signal ptr_deref_5137_store_0_req_0 : boolean;
  signal type_cast_3008_inst_ack_1 : boolean;
  signal ptr_deref_5137_store_0_ack_0 : boolean;
  signal ptr_deref_5137_store_0_req_1 : boolean;
  signal phi_stmt_3005_req_0 : boolean;
  signal ptr_deref_5137_store_0_ack_1 : boolean;
  signal type_cast_5145_inst_req_0 : boolean;
  signal type_cast_5145_inst_ack_0 : boolean;
  signal type_cast_5145_inst_req_1 : boolean;
  signal type_cast_5145_inst_ack_1 : boolean;
  signal if_stmt_5160_branch_req_0 : boolean;
  signal if_stmt_5160_branch_ack_1 : boolean;
  signal if_stmt_5160_branch_ack_0 : boolean;
  signal type_cast_5184_inst_req_0 : boolean;
  signal type_cast_5184_inst_ack_0 : boolean;
  signal type_cast_5184_inst_req_1 : boolean;
  signal type_cast_5184_inst_ack_1 : boolean;
  signal type_cast_2986_inst_req_0 : boolean;
  signal LOAD_col_high_5187_load_0_req_0 : boolean;
  signal LOAD_col_high_5187_load_0_ack_0 : boolean;
  signal LOAD_col_high_5187_load_0_req_1 : boolean;
  signal LOAD_col_high_5187_load_0_ack_1 : boolean;
  signal type_cast_5191_inst_req_0 : boolean;
  signal type_cast_5191_inst_ack_0 : boolean;
  signal type_cast_5191_inst_req_1 : boolean;
  signal type_cast_5191_inst_ack_1 : boolean;
  signal type_cast_5205_inst_req_0 : boolean;
  signal type_cast_5205_inst_ack_0 : boolean;
  signal type_cast_5205_inst_req_1 : boolean;
  signal type_cast_5205_inst_ack_1 : boolean;
  signal type_cast_5221_inst_req_0 : boolean;
  signal type_cast_5221_inst_ack_0 : boolean;
  signal type_cast_5221_inst_req_1 : boolean;
  signal phi_stmt_1307_req_1 : boolean;
  signal phi_stmt_1307_ack_0 : boolean;
  signal phi_stmt_1313_ack_0 : boolean;
  signal phi_stmt_1319_ack_0 : boolean;
  signal type_cast_1332_inst_req_0 : boolean;
  signal type_cast_1332_inst_ack_0 : boolean;
  signal type_cast_1332_inst_req_1 : boolean;
  signal type_cast_1332_inst_ack_1 : boolean;
  signal phi_stmt_1329_req_0 : boolean;
  signal type_cast_1336_inst_req_0 : boolean;
  signal type_cast_1336_inst_ack_0 : boolean;
  signal type_cast_1336_inst_req_1 : boolean;
  signal type_cast_1336_inst_ack_1 : boolean;
  signal phi_stmt_1333_req_0 : boolean;
  signal phi_stmt_1329_ack_0 : boolean;
  signal phi_stmt_1333_ack_0 : boolean;
  signal type_cast_1469_inst_req_0 : boolean;
  signal type_cast_1469_inst_ack_0 : boolean;
  signal type_cast_1469_inst_req_1 : boolean;
  signal type_cast_1469_inst_ack_1 : boolean;
  signal phi_stmt_1464_req_1 : boolean;
  signal type_cast_1476_inst_req_0 : boolean;
  signal type_cast_1476_inst_ack_0 : boolean;
  signal type_cast_1476_inst_req_1 : boolean;
  signal type_cast_1476_inst_ack_1 : boolean;
  signal phi_stmt_1470_req_1 : boolean;
  signal type_cast_1483_inst_req_0 : boolean;
  signal type_cast_1483_inst_ack_0 : boolean;
  signal type_cast_1483_inst_req_1 : boolean;
  signal type_cast_1483_inst_ack_1 : boolean;
  signal phi_stmt_1477_req_1 : boolean;
  signal type_cast_1467_inst_req_0 : boolean;
  signal type_cast_1467_inst_ack_0 : boolean;
  signal type_cast_1467_inst_req_1 : boolean;
  signal type_cast_1467_inst_ack_1 : boolean;
  signal phi_stmt_1464_req_0 : boolean;
  signal phi_stmt_1470_req_0 : boolean;
  signal phi_stmt_1477_req_0 : boolean;
  signal phi_stmt_1464_ack_0 : boolean;
  signal phi_stmt_1470_ack_0 : boolean;
  signal phi_stmt_1477_ack_0 : boolean;
  signal phi_stmt_1869_req_1 : boolean;
  signal type_cast_1868_inst_req_0 : boolean;
  signal type_cast_1868_inst_ack_0 : boolean;
  signal phi_stmt_3147_req_0 : boolean;
  signal type_cast_1868_inst_req_1 : boolean;
  signal type_cast_1868_inst_ack_1 : boolean;
  signal phi_stmt_2990_req_1 : boolean;
  signal phi_stmt_1863_req_1 : boolean;
  signal type_cast_2995_inst_ack_1 : boolean;
  signal type_cast_2995_inst_req_1 : boolean;
  signal type_cast_3150_inst_ack_1 : boolean;
  signal type_cast_1862_inst_req_0 : boolean;
  signal type_cast_1862_inst_ack_0 : boolean;
  signal type_cast_3150_inst_req_1 : boolean;
  signal type_cast_1862_inst_req_1 : boolean;
  signal type_cast_1862_inst_ack_1 : boolean;
  signal type_cast_2995_inst_ack_0 : boolean;
  signal phi_stmt_1857_req_1 : boolean;
  signal type_cast_2995_inst_req_0 : boolean;
  signal type_cast_1872_inst_req_0 : boolean;
  signal type_cast_1872_inst_ack_0 : boolean;
  signal type_cast_1872_inst_req_1 : boolean;
  signal type_cast_1872_inst_ack_1 : boolean;
  signal phi_stmt_1869_req_0 : boolean;
  signal type_cast_3150_inst_ack_0 : boolean;
  signal type_cast_1866_inst_req_0 : boolean;
  signal type_cast_1866_inst_ack_0 : boolean;
  signal type_cast_1866_inst_req_1 : boolean;
  signal type_cast_3008_inst_req_1 : boolean;
  signal type_cast_1866_inst_ack_1 : boolean;
  signal phi_stmt_1863_req_0 : boolean;
  signal type_cast_3150_inst_req_0 : boolean;
  signal type_cast_1860_inst_req_0 : boolean;
  signal type_cast_1860_inst_ack_0 : boolean;
  signal type_cast_1860_inst_req_1 : boolean;
  signal type_cast_1860_inst_ack_1 : boolean;
  signal phi_stmt_1857_req_0 : boolean;
  signal type_cast_3008_inst_ack_0 : boolean;
  signal phi_stmt_1857_ack_0 : boolean;
  signal phi_stmt_1863_ack_0 : boolean;
  signal phi_stmt_1869_ack_0 : boolean;
  signal type_cast_1886_inst_req_0 : boolean;
  signal type_cast_1886_inst_ack_0 : boolean;
  signal type_cast_3008_inst_req_0 : boolean;
  signal type_cast_1886_inst_req_1 : boolean;
  signal type_cast_1886_inst_ack_1 : boolean;
  signal phi_stmt_1883_req_0 : boolean;
  signal phi_stmt_3153_ack_0 : boolean;
  signal phi_stmt_3147_ack_0 : boolean;
  signal type_cast_1882_inst_req_0 : boolean;
  signal type_cast_1882_inst_ack_0 : boolean;
  signal type_cast_1882_inst_req_1 : boolean;
  signal type_cast_1882_inst_ack_1 : boolean;
  signal phi_stmt_1879_req_0 : boolean;
  signal phi_stmt_1879_ack_0 : boolean;
  signal phi_stmt_1883_ack_0 : boolean;
  signal phi_stmt_2983_req_1 : boolean;
  signal phi_stmt_3140_ack_0 : boolean;
  signal type_cast_2030_inst_req_0 : boolean;
  signal type_cast_2030_inst_ack_0 : boolean;
  signal type_cast_2030_inst_req_1 : boolean;
  signal type_cast_2030_inst_ack_1 : boolean;
  signal phi_stmt_2027_req_0 : boolean;
  signal type_cast_2017_inst_req_0 : boolean;
  signal type_cast_2017_inst_ack_0 : boolean;
  signal type_cast_2017_inst_req_1 : boolean;
  signal type_cast_2017_inst_ack_1 : boolean;
  signal phi_stmt_2014_req_0 : boolean;
  signal phi_stmt_3140_req_0 : boolean;
  signal type_cast_2026_inst_req_0 : boolean;
  signal type_cast_2026_inst_ack_0 : boolean;
  signal type_cast_2026_inst_req_1 : boolean;
  signal type_cast_2026_inst_ack_1 : boolean;
  signal phi_stmt_2021_req_1 : boolean;
  signal phi_stmt_3140_req_1 : boolean;
  signal type_cast_3146_inst_ack_1 : boolean;
  signal phi_stmt_2027_req_1 : boolean;
  signal type_cast_3146_inst_req_1 : boolean;
  signal phi_stmt_2014_req_1 : boolean;
  signal type_cast_2024_inst_req_0 : boolean;
  signal phi_stmt_3153_req_0 : boolean;
  signal type_cast_2024_inst_ack_0 : boolean;
  signal phi_stmt_2996_ack_0 : boolean;
  signal type_cast_2024_inst_req_1 : boolean;
  signal phi_stmt_2990_ack_0 : boolean;
  signal type_cast_2024_inst_ack_1 : boolean;
  signal phi_stmt_2021_req_0 : boolean;
  signal type_cast_3156_inst_ack_1 : boolean;
  signal phi_stmt_2983_ack_0 : boolean;
  signal type_cast_3156_inst_req_1 : boolean;
  signal phi_stmt_2014_ack_0 : boolean;
  signal phi_stmt_2021_ack_0 : boolean;
  signal phi_stmt_2027_ack_0 : boolean;
  signal phi_stmt_2983_req_0 : boolean;
  signal phi_stmt_2996_req_0 : boolean;
  signal type_cast_4877_inst_req_0 : boolean;
  signal phi_stmt_2996_req_1 : boolean;
  signal type_cast_3001_inst_ack_1 : boolean;
  signal type_cast_2999_inst_ack_1 : boolean;
  signal phi_stmt_3147_req_1 : boolean;
  signal type_cast_2999_inst_req_1 : boolean;
  signal type_cast_3152_inst_ack_1 : boolean;
  signal type_cast_3152_inst_req_1 : boolean;
  signal type_cast_2999_inst_ack_0 : boolean;
  signal type_cast_2999_inst_req_0 : boolean;
  signal phi_stmt_3153_req_1 : boolean;
  signal type_cast_3001_inst_req_1 : boolean;
  signal type_cast_3001_inst_ack_0 : boolean;
  signal type_cast_2986_inst_ack_1 : boolean;
  signal type_cast_3001_inst_req_0 : boolean;
  signal type_cast_2986_inst_req_1 : boolean;
  signal type_cast_3146_inst_ack_0 : boolean;
  signal phi_stmt_2990_req_0 : boolean;
  signal type_cast_3156_inst_ack_0 : boolean;
  signal type_cast_3152_inst_ack_0 : boolean;
  signal type_cast_3146_inst_req_0 : boolean;
  signal phi_stmt_2420_req_1 : boolean;
  signal type_cast_3152_inst_req_0 : boolean;
  signal type_cast_2432_inst_req_0 : boolean;
  signal type_cast_3156_inst_req_0 : boolean;
  signal type_cast_2432_inst_ack_0 : boolean;
  signal type_cast_2993_inst_ack_1 : boolean;
  signal type_cast_2432_inst_req_1 : boolean;
  signal type_cast_2993_inst_req_1 : boolean;
  signal type_cast_2432_inst_ack_1 : boolean;
  signal phi_stmt_2427_req_1 : boolean;
  signal type_cast_2986_inst_ack_0 : boolean;
  signal type_cast_2438_inst_req_0 : boolean;
  signal type_cast_2438_inst_ack_0 : boolean;
  signal type_cast_2438_inst_req_1 : boolean;
  signal type_cast_2438_inst_ack_1 : boolean;
  signal phi_stmt_2433_req_1 : boolean;
  signal type_cast_2993_inst_ack_0 : boolean;
  signal type_cast_2423_inst_req_0 : boolean;
  signal type_cast_2423_inst_ack_0 : boolean;
  signal type_cast_2993_inst_req_0 : boolean;
  signal type_cast_2423_inst_req_1 : boolean;
  signal type_cast_2423_inst_ack_1 : boolean;
  signal phi_stmt_2420_req_0 : boolean;
  signal type_cast_2430_inst_req_0 : boolean;
  signal type_cast_2430_inst_ack_0 : boolean;
  signal type_cast_2430_inst_req_1 : boolean;
  signal type_cast_2430_inst_ack_1 : boolean;
  signal phi_stmt_2427_req_0 : boolean;
  signal type_cast_2436_inst_req_0 : boolean;
  signal type_cast_2436_inst_ack_0 : boolean;
  signal type_cast_2436_inst_req_1 : boolean;
  signal type_cast_2436_inst_ack_1 : boolean;
  signal phi_stmt_2433_req_0 : boolean;
  signal phi_stmt_2420_ack_0 : boolean;
  signal phi_stmt_2427_ack_0 : boolean;
  signal phi_stmt_2433_ack_0 : boolean;
  signal type_cast_5263_inst_req_0 : boolean;
  signal type_cast_2445_inst_req_0 : boolean;
  signal type_cast_5263_inst_ack_0 : boolean;
  signal type_cast_2445_inst_ack_0 : boolean;
  signal type_cast_2445_inst_req_1 : boolean;
  signal type_cast_2445_inst_ack_1 : boolean;
  signal phi_stmt_2442_req_0 : boolean;
  signal type_cast_2449_inst_req_0 : boolean;
  signal type_cast_2449_inst_ack_0 : boolean;
  signal type_cast_2449_inst_req_1 : boolean;
  signal type_cast_2449_inst_ack_1 : boolean;
  signal phi_stmt_2446_req_0 : boolean;
  signal type_cast_2453_inst_req_0 : boolean;
  signal type_cast_2453_inst_ack_0 : boolean;
  signal type_cast_2453_inst_req_1 : boolean;
  signal type_cast_2453_inst_ack_1 : boolean;
  signal phi_stmt_2450_req_0 : boolean;
  signal phi_stmt_2442_ack_0 : boolean;
  signal phi_stmt_2446_ack_0 : boolean;
  signal phi_stmt_2450_ack_0 : boolean;
  signal type_cast_2597_inst_req_0 : boolean;
  signal type_cast_2597_inst_ack_0 : boolean;
  signal type_cast_2597_inst_req_1 : boolean;
  signal type_cast_2597_inst_ack_1 : boolean;
  signal phi_stmt_2591_req_1 : boolean;
  signal type_cast_2603_inst_req_0 : boolean;
  signal type_cast_2603_inst_ack_0 : boolean;
  signal type_cast_2603_inst_req_1 : boolean;
  signal type_cast_2603_inst_ack_1 : boolean;
  signal phi_stmt_2598_req_1 : boolean;
  signal type_cast_5263_inst_req_1 : boolean;
  signal type_cast_2609_inst_req_0 : boolean;
  signal type_cast_2609_inst_ack_0 : boolean;
  signal type_cast_2609_inst_req_1 : boolean;
  signal type_cast_2609_inst_ack_1 : boolean;
  signal phi_stmt_2604_req_1 : boolean;
  signal type_cast_5265_inst_req_0 : boolean;
  signal phi_stmt_2591_req_0 : boolean;
  signal type_cast_2601_inst_req_0 : boolean;
  signal type_cast_5263_inst_ack_1 : boolean;
  signal type_cast_2601_inst_ack_0 : boolean;
  signal type_cast_2601_inst_req_1 : boolean;
  signal type_cast_2601_inst_ack_1 : boolean;
  signal phi_stmt_2598_req_0 : boolean;
  signal type_cast_2607_inst_req_0 : boolean;
  signal type_cast_2607_inst_ack_0 : boolean;
  signal type_cast_2607_inst_req_1 : boolean;
  signal type_cast_2607_inst_ack_1 : boolean;
  signal phi_stmt_2604_req_0 : boolean;
  signal phi_stmt_2591_ack_0 : boolean;
  signal phi_stmt_2598_ack_0 : boolean;
  signal phi_stmt_2604_ack_0 : boolean;
  signal phi_stmt_3558_req_1 : boolean;
  signal type_cast_3570_inst_req_0 : boolean;
  signal type_cast_3570_inst_ack_0 : boolean;
  signal type_cast_3570_inst_req_1 : boolean;
  signal type_cast_3570_inst_ack_1 : boolean;
  signal phi_stmt_3565_req_1 : boolean;
  signal type_cast_3574_inst_req_0 : boolean;
  signal type_cast_3574_inst_ack_0 : boolean;
  signal type_cast_3574_inst_req_1 : boolean;
  signal type_cast_3574_inst_ack_1 : boolean;
  signal phi_stmt_3571_req_0 : boolean;
  signal type_cast_3561_inst_req_0 : boolean;
  signal type_cast_3561_inst_ack_0 : boolean;
  signal type_cast_3561_inst_req_1 : boolean;
  signal type_cast_3561_inst_ack_1 : boolean;
  signal phi_stmt_3558_req_0 : boolean;
  signal type_cast_3568_inst_req_0 : boolean;
  signal type_cast_3568_inst_ack_0 : boolean;
  signal type_cast_3568_inst_req_1 : boolean;
  signal type_cast_3568_inst_ack_1 : boolean;
  signal phi_stmt_3565_req_0 : boolean;
  signal type_cast_3576_inst_req_0 : boolean;
  signal type_cast_3576_inst_ack_0 : boolean;
  signal type_cast_3576_inst_req_1 : boolean;
  signal type_cast_3576_inst_ack_1 : boolean;
  signal phi_stmt_3571_req_1 : boolean;
  signal phi_stmt_3558_ack_0 : boolean;
  signal phi_stmt_3565_ack_0 : boolean;
  signal phi_stmt_3571_ack_0 : boolean;
  signal type_cast_3583_inst_req_0 : boolean;
  signal type_cast_3583_inst_ack_0 : boolean;
  signal type_cast_3583_inst_req_1 : boolean;
  signal type_cast_3583_inst_ack_1 : boolean;
  signal phi_stmt_3580_req_0 : boolean;
  signal type_cast_3587_inst_req_0 : boolean;
  signal type_cast_3587_inst_ack_0 : boolean;
  signal type_cast_3587_inst_req_1 : boolean;
  signal type_cast_3587_inst_ack_1 : boolean;
  signal phi_stmt_3584_req_0 : boolean;
  signal type_cast_3591_inst_req_0 : boolean;
  signal type_cast_3591_inst_ack_0 : boolean;
  signal type_cast_3591_inst_req_1 : boolean;
  signal type_cast_3591_inst_ack_1 : boolean;
  signal phi_stmt_3588_req_0 : boolean;
  signal phi_stmt_3580_ack_0 : boolean;
  signal phi_stmt_3584_ack_0 : boolean;
  signal phi_stmt_3588_ack_0 : boolean;
  signal type_cast_3732_inst_req_0 : boolean;
  signal type_cast_3732_inst_ack_0 : boolean;
  signal type_cast_3732_inst_req_1 : boolean;
  signal type_cast_3732_inst_ack_1 : boolean;
  signal phi_stmt_3729_req_0 : boolean;
  signal type_cast_3739_inst_req_0 : boolean;
  signal type_cast_3739_inst_ack_0 : boolean;
  signal type_cast_3739_inst_req_1 : boolean;
  signal type_cast_3739_inst_ack_1 : boolean;
  signal phi_stmt_3736_req_0 : boolean;
  signal type_cast_3747_inst_req_0 : boolean;
  signal type_cast_3747_inst_ack_0 : boolean;
  signal type_cast_3747_inst_req_1 : boolean;
  signal type_cast_3747_inst_ack_1 : boolean;
  signal phi_stmt_3742_req_1 : boolean;
  signal phi_stmt_3729_req_1 : boolean;
  signal type_cast_3741_inst_req_0 : boolean;
  signal type_cast_3741_inst_ack_0 : boolean;
  signal type_cast_3741_inst_req_1 : boolean;
  signal type_cast_3741_inst_ack_1 : boolean;
  signal phi_stmt_3736_req_1 : boolean;
  signal type_cast_3745_inst_req_0 : boolean;
  signal type_cast_3745_inst_ack_0 : boolean;
  signal type_cast_3745_inst_req_1 : boolean;
  signal type_cast_3745_inst_ack_1 : boolean;
  signal phi_stmt_3742_req_0 : boolean;
  signal phi_stmt_3729_ack_0 : boolean;
  signal phi_stmt_3736_ack_0 : boolean;
  signal phi_stmt_3742_ack_0 : boolean;
  signal phi_stmt_4880_req_1 : boolean;
  signal type_cast_4885_inst_ack_1 : boolean;
  signal type_cast_5250_inst_ack_0 : boolean;
  signal type_cast_5250_inst_req_0 : boolean;
  signal type_cast_4885_inst_req_1 : boolean;
  signal type_cast_4885_inst_ack_0 : boolean;
  signal type_cast_4885_inst_req_0 : boolean;
  signal phi_stmt_4133_req_1 : boolean;
  signal type_cast_4145_inst_req_0 : boolean;
  signal type_cast_4145_inst_ack_0 : boolean;
  signal type_cast_4145_inst_req_1 : boolean;
  signal type_cast_4145_inst_ack_1 : boolean;
  signal phi_stmt_4140_req_1 : boolean;
  signal type_cast_4151_inst_req_0 : boolean;
  signal type_cast_4151_inst_ack_0 : boolean;
  signal type_cast_4151_inst_req_1 : boolean;
  signal type_cast_4151_inst_ack_1 : boolean;
  signal phi_stmt_4146_req_1 : boolean;
  signal type_cast_4136_inst_req_0 : boolean;
  signal type_cast_4136_inst_ack_0 : boolean;
  signal type_cast_4136_inst_req_1 : boolean;
  signal type_cast_4136_inst_ack_1 : boolean;
  signal phi_stmt_4133_req_0 : boolean;
  signal phi_stmt_5254_req_0 : boolean;
  signal type_cast_5257_inst_ack_1 : boolean;
  signal type_cast_4143_inst_req_0 : boolean;
  signal phi_stmt_5254_req_1 : boolean;
  signal type_cast_4143_inst_ack_0 : boolean;
  signal type_cast_4143_inst_req_1 : boolean;
  signal type_cast_4143_inst_ack_1 : boolean;
  signal phi_stmt_4140_req_0 : boolean;
  signal type_cast_5259_inst_ack_1 : boolean;
  signal type_cast_5257_inst_req_1 : boolean;
  signal type_cast_4149_inst_req_0 : boolean;
  signal type_cast_5259_inst_req_1 : boolean;
  signal type_cast_4149_inst_ack_0 : boolean;
  signal type_cast_4149_inst_req_1 : boolean;
  signal type_cast_4149_inst_ack_1 : boolean;
  signal phi_stmt_4146_req_0 : boolean;
  signal phi_stmt_4133_ack_0 : boolean;
  signal phi_stmt_5260_req_0 : boolean;
  signal phi_stmt_4140_ack_0 : boolean;
  signal phi_stmt_4146_ack_0 : boolean;
  signal phi_stmt_4880_ack_0 : boolean;
  signal type_cast_5257_inst_ack_0 : boolean;
  signal type_cast_5257_inst_req_0 : boolean;
  signal type_cast_4158_inst_req_0 : boolean;
  signal type_cast_4158_inst_ack_0 : boolean;
  signal type_cast_4158_inst_req_1 : boolean;
  signal type_cast_4158_inst_ack_1 : boolean;
  signal phi_stmt_5260_req_1 : boolean;
  signal phi_stmt_4155_req_0 : boolean;
  signal phi_stmt_4874_ack_0 : boolean;
  signal phi_stmt_4874_req_0 : boolean;
  signal type_cast_4877_inst_ack_1 : boolean;
  signal type_cast_4162_inst_req_0 : boolean;
  signal type_cast_4162_inst_ack_0 : boolean;
  signal type_cast_5259_inst_ack_0 : boolean;
  signal type_cast_4162_inst_req_1 : boolean;
  signal type_cast_4162_inst_ack_1 : boolean;
  signal type_cast_4877_inst_req_1 : boolean;
  signal phi_stmt_4159_req_0 : boolean;
  signal type_cast_5259_inst_req_0 : boolean;
  signal phi_stmt_4155_ack_0 : boolean;
  signal phi_stmt_4159_ack_0 : boolean;
  signal phi_stmt_4867_ack_0 : boolean;
  signal type_cast_4302_inst_req_0 : boolean;
  signal type_cast_4302_inst_ack_0 : boolean;
  signal type_cast_4302_inst_req_1 : boolean;
  signal type_cast_4302_inst_ack_1 : boolean;
  signal type_cast_5265_inst_ack_1 : boolean;
  signal phi_stmt_4296_req_1 : boolean;
  signal type_cast_4308_inst_req_0 : boolean;
  signal type_cast_4308_inst_ack_0 : boolean;
  signal type_cast_4308_inst_req_1 : boolean;
  signal type_cast_4308_inst_ack_1 : boolean;
  signal phi_stmt_4303_req_1 : boolean;
  signal type_cast_4315_inst_req_0 : boolean;
  signal type_cast_4315_inst_ack_0 : boolean;
  signal type_cast_4315_inst_req_1 : boolean;
  signal type_cast_4315_inst_ack_1 : boolean;
  signal phi_stmt_4309_req_1 : boolean;
  signal phi_stmt_4296_req_0 : boolean;
  signal phi_stmt_5247_req_0 : boolean;
  signal type_cast_4306_inst_req_0 : boolean;
  signal type_cast_4306_inst_ack_0 : boolean;
  signal type_cast_4306_inst_req_1 : boolean;
  signal type_cast_4306_inst_ack_1 : boolean;
  signal phi_stmt_4303_req_0 : boolean;
  signal phi_stmt_4309_req_0 : boolean;
  signal type_cast_5250_inst_ack_1 : boolean;
  signal type_cast_5265_inst_req_1 : boolean;
  signal phi_stmt_4296_ack_0 : boolean;
  signal phi_stmt_4303_ack_0 : boolean;
  signal phi_stmt_4309_ack_0 : boolean;
  signal phi_stmt_4867_req_0 : boolean;
  signal phi_stmt_5247_req_1 : boolean;
  signal type_cast_4877_inst_ack_0 : boolean;
  signal type_cast_5250_inst_req_1 : boolean;
  signal type_cast_5265_inst_ack_0 : boolean;
  signal type_cast_4706_inst_req_0 : boolean;
  signal type_cast_4706_inst_ack_0 : boolean;
  signal type_cast_4706_inst_req_1 : boolean;
  signal type_cast_4706_inst_ack_1 : boolean;
  signal phi_stmt_4703_req_0 : boolean;
  signal type_cast_4702_inst_req_0 : boolean;
  signal type_cast_4702_inst_ack_0 : boolean;
  signal type_cast_4702_inst_req_1 : boolean;
  signal type_cast_4702_inst_ack_1 : boolean;
  signal phi_stmt_4697_req_1 : boolean;
  signal phi_stmt_4690_req_0 : boolean;
  signal type_cast_4708_inst_req_0 : boolean;
  signal type_cast_4708_inst_ack_0 : boolean;
  signal type_cast_4708_inst_req_1 : boolean;
  signal type_cast_4708_inst_ack_1 : boolean;
  signal phi_stmt_4703_req_1 : boolean;
  signal type_cast_4700_inst_req_0 : boolean;
  signal type_cast_4700_inst_ack_0 : boolean;
  signal type_cast_4700_inst_req_1 : boolean;
  signal type_cast_4700_inst_ack_1 : boolean;
  signal phi_stmt_4697_req_0 : boolean;
  signal type_cast_4696_inst_req_0 : boolean;
  signal type_cast_4696_inst_ack_0 : boolean;
  signal type_cast_4696_inst_req_1 : boolean;
  signal type_cast_4696_inst_ack_1 : boolean;
  signal phi_stmt_4690_req_1 : boolean;
  signal phi_stmt_4690_ack_0 : boolean;
  signal phi_stmt_4697_ack_0 : boolean;
  signal phi_stmt_4703_ack_0 : boolean;
  signal type_cast_4719_inst_req_0 : boolean;
  signal type_cast_4719_inst_ack_0 : boolean;
  signal type_cast_4719_inst_req_1 : boolean;
  signal type_cast_4719_inst_ack_1 : boolean;
  signal phi_stmt_4716_req_0 : boolean;
  signal type_cast_4715_inst_req_0 : boolean;
  signal type_cast_4715_inst_ack_0 : boolean;
  signal type_cast_4715_inst_req_1 : boolean;
  signal type_cast_4715_inst_ack_1 : boolean;
  signal phi_stmt_4712_req_0 : boolean;
  signal type_cast_4723_inst_req_0 : boolean;
  signal type_cast_4723_inst_ack_0 : boolean;
  signal type_cast_4723_inst_req_1 : boolean;
  signal type_cast_4723_inst_ack_1 : boolean;
  signal phi_stmt_4720_req_0 : boolean;
  signal phi_stmt_4712_ack_0 : boolean;
  signal phi_stmt_4716_ack_0 : boolean;
  signal phi_stmt_4720_ack_0 : boolean;
  signal type_cast_4879_inst_req_0 : boolean;
  signal type_cast_4879_inst_ack_0 : boolean;
  signal type_cast_4879_inst_req_1 : boolean;
  signal type_cast_4879_inst_ack_1 : boolean;
  signal phi_stmt_4874_req_1 : boolean;
  signal type_cast_4883_inst_req_0 : boolean;
  signal type_cast_4883_inst_ack_0 : boolean;
  signal type_cast_4883_inst_req_1 : boolean;
  signal type_cast_4883_inst_ack_1 : boolean;
  signal phi_stmt_4880_req_0 : boolean;
  signal type_cast_4873_inst_req_0 : boolean;
  signal type_cast_4873_inst_ack_0 : boolean;
  signal type_cast_4873_inst_req_1 : boolean;
  signal type_cast_4873_inst_ack_1 : boolean;
  signal phi_stmt_4867_req_1 : boolean;
  signal phi_stmt_5247_ack_0 : boolean;
  signal phi_stmt_5254_ack_0 : boolean;
  signal phi_stmt_5260_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_CP_2152_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_2152_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_CP_2152_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_2152_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_CP_2152: Block -- control-path 
    signal zeropad3D_CP_2152_elements: BooleanArray(1233 downto 0);
    -- 
  begin -- 
    zeropad3D_CP_2152_elements(0) <= zeropad3D_CP_2152_start;
    zeropad3D_CP_2152_symbol <= zeropad3D_CP_2152_elements(779);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	15 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	18 
    -- CP-element group 0: 	19 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	26 
    -- CP-element group 0: 	27 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	31 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	34 
    -- CP-element group 0:  members (104) 
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773__entry__
      -- CP-element group 0: 	 branch_block_stmt_714/branch_block_stmt_714__entry__
      -- CP-element group 0: 	 branch_block_stmt_714/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Update/ccr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/word_access_complete/word_0/cr
      -- 
    crr_2608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => call_stmt_716_call_req_0); -- 
    ccr_2613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => call_stmt_716_call_req_1); -- 
    cr_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => ptr_deref_727_load_0_req_1); -- 
    cr_2677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => type_cast_731_inst_req_1); -- 
    cr_2710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => STORE_row_high_733_store_0_req_1); -- 
    cr_2755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => ptr_deref_746_load_0_req_1); -- 
    cr_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => type_cast_750_inst_req_1); -- 
    cr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => STORE_col_high_752_store_0_req_1); -- 
    cr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => ptr_deref_765_load_0_req_1); -- 
    cr_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => type_cast_769_inst_req_1); -- 
    cr_2904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => STORE_depth_high_771_store_0_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	823 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	784 
    -- CP-element group 1: 	785 
    -- CP-element group 1: 	787 
    -- CP-element group 1: 	788 
    -- CP-element group 1: 	790 
    -- CP-element group 1: 	791 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_714/merge_stmt_1306__exit__
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/$entry
      -- 
    cr_11022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1), ack => type_cast_905_inst_req_1); -- 
    rr_11017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1), ack => type_cast_905_inst_req_0); -- 
    cr_11045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1), ack => type_cast_912_inst_req_1); -- 
    rr_11040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1), ack => type_cast_912_inst_req_0); -- 
    cr_11068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1), ack => type_cast_919_inst_req_1); -- 
    rr_11063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1), ack => type_cast_919_inst_req_0); -- 
    zeropad3D_CP_2152_elements(1) <= zeropad3D_CP_2152_elements(823);
    -- CP-element group 2:  merge  fork  transition  place  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	879 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	834 
    -- CP-element group 2: 	835 
    -- CP-element group 2: 	837 
    -- CP-element group 2: 	838 
    -- CP-element group 2: 	840 
    -- CP-element group 2: 	841 
    -- CP-element group 2:  members (27) 
      -- CP-element group 2: 	 branch_block_stmt_714/merge_stmt_1856__exit__
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1469/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1469/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1469/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1469/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1469/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1469/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/type_cast_1476/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/type_cast_1476/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/type_cast_1476/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/type_cast_1476/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/type_cast_1476/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/type_cast_1476/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/type_cast_1483/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/type_cast_1483/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/type_cast_1483/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/type_cast_1483/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/type_cast_1483/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/type_cast_1483/SplitProtocol/Update/cr
      -- 
    rr_11387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(2), ack => type_cast_1469_inst_req_0); -- 
    cr_11392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(2), ack => type_cast_1469_inst_req_1); -- 
    rr_11410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(2), ack => type_cast_1476_inst_req_0); -- 
    cr_11415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(2), ack => type_cast_1476_inst_req_1); -- 
    rr_11433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(2), ack => type_cast_1483_inst_req_0); -- 
    cr_11438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(2), ack => type_cast_1483_inst_req_1); -- 
    zeropad3D_CP_2152_elements(2) <= zeropad3D_CP_2152_elements(879);
    -- CP-element group 3:  merge  fork  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	935 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	890 
    -- CP-element group 3: 	891 
    -- CP-element group 3: 	893 
    -- CP-element group 3: 	894 
    -- CP-element group 3: 	896 
    -- CP-element group 3: 	897 
    -- CP-element group 3:  members (27) 
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460
      -- CP-element group 3: 	 branch_block_stmt_714/merge_stmt_2419__exit__
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/type_cast_2030/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/type_cast_2030/SplitProtocol/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/type_cast_2030/SplitProtocol/Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/type_cast_2030/SplitProtocol/Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/type_cast_2030/SplitProtocol/Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/type_cast_2030/SplitProtocol/Update/cr
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Update/cr
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2026/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2026/SplitProtocol/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2026/SplitProtocol/Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2026/SplitProtocol/Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2026/SplitProtocol/Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2026/SplitProtocol/Update/cr
      -- 
    rr_11799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(3), ack => type_cast_2030_inst_req_0); -- 
    cr_11804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(3), ack => type_cast_2030_inst_req_1); -- 
    rr_11822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(3), ack => type_cast_2017_inst_req_0); -- 
    cr_11827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(3), ack => type_cast_2017_inst_req_1); -- 
    rr_11845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(3), ack => type_cast_2026_inst_req_0); -- 
    cr_11850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(3), ack => type_cast_2026_inst_req_1); -- 
    zeropad3D_CP_2152_elements(3) <= zeropad3D_CP_2152_elements(935);
    -- CP-element group 4:  merge  fork  transition  place  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	997 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	950 
    -- CP-element group 4: 	951 
    -- CP-element group 4: 	953 
    -- CP-element group 4: 	954 
    -- CP-element group 4: 	956 
    -- CP-element group 4: 	957 
    -- CP-element group 4:  members (27) 
      -- CP-element group 4: 	 branch_block_stmt_714/merge_stmt_2982__exit__
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/type_cast_2597/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/type_cast_2597/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/type_cast_2597/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/type_cast_2597/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/type_cast_2597/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/type_cast_2597/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2603/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2603/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2603/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2603/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2603/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2603/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2609/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2609/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2609/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2609/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2609/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2609/SplitProtocol/Update/cr
      -- 
    rr_12235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(4), ack => type_cast_2597_inst_req_0); -- 
    cr_12240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(4), ack => type_cast_2597_inst_req_1); -- 
    rr_12258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(4), ack => type_cast_2603_inst_req_0); -- 
    cr_12263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(4), ack => type_cast_2603_inst_req_1); -- 
    rr_12281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(4), ack => type_cast_2609_inst_req_0); -- 
    cr_12286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(4), ack => type_cast_2609_inst_req_1); -- 
    zeropad3D_CP_2152_elements(4) <= zeropad3D_CP_2152_elements(997);
    -- CP-element group 5:  merge  fork  transition  place  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1053 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	1008 
    -- CP-element group 5: 	1009 
    -- CP-element group 5: 	1011 
    -- CP-element group 5: 	1012 
    -- CP-element group 5: 	1014 
    -- CP-element group 5: 	1015 
    -- CP-element group 5:  members (27) 
      -- CP-element group 5: 	 branch_block_stmt_714/merge_stmt_3557__exit__
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/type_cast_3156/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/type_cast_3146/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3150/SplitProtocol/Update/cr
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3150/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3150/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/type_cast_3146/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/type_cast_3146/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/type_cast_3156/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3150/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3150/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3150/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/type_cast_3146/SplitProtocol/Update/cr
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/type_cast_3156/SplitProtocol/Update/cr
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/type_cast_3156/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/type_cast_3146/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/type_cast_3146/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/type_cast_3156/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/type_cast_3156/SplitProtocol/Sample/$entry
      -- 
    cr_12690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(5), ack => type_cast_3150_inst_req_1); -- 
    rr_12685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(5), ack => type_cast_3150_inst_req_0); -- 
    cr_12713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(5), ack => type_cast_3146_inst_req_1); -- 
    cr_12667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(5), ack => type_cast_3156_inst_req_1); -- 
    rr_12708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(5), ack => type_cast_3146_inst_req_0); -- 
    rr_12662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(5), ack => type_cast_3156_inst_req_0); -- 
    zeropad3D_CP_2152_elements(5) <= zeropad3D_CP_2152_elements(1053);
    -- CP-element group 6:  merge  fork  transition  place  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1115 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	1068 
    -- CP-element group 6: 	1069 
    -- CP-element group 6: 	1071 
    -- CP-element group 6: 	1072 
    -- CP-element group 6: 	1074 
    -- CP-element group 6: 	1075 
    -- CP-element group 6:  members (27) 
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122
      -- CP-element group 6: 	 branch_block_stmt_714/merge_stmt_4132__exit__
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/type_cast_3732/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/type_cast_3732/SplitProtocol/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/type_cast_3732/SplitProtocol/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/type_cast_3732/SplitProtocol/Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/type_cast_3732/SplitProtocol/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/type_cast_3732/SplitProtocol/Update/cr
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3739/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3739/SplitProtocol/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3739/SplitProtocol/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3739/SplitProtocol/Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3739/SplitProtocol/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3739/SplitProtocol/Update/cr
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3747/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3747/SplitProtocol/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3747/SplitProtocol/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3747/SplitProtocol/Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3747/SplitProtocol/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3747/SplitProtocol/Update/cr
      -- 
    rr_13098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(6), ack => type_cast_3732_inst_req_0); -- 
    cr_13103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(6), ack => type_cast_3732_inst_req_1); -- 
    rr_13121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(6), ack => type_cast_3739_inst_req_0); -- 
    cr_13126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(6), ack => type_cast_3739_inst_req_1); -- 
    rr_13144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(6), ack => type_cast_3747_inst_req_0); -- 
    cr_13149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(6), ack => type_cast_3747_inst_req_1); -- 
    zeropad3D_CP_2152_elements(6) <= zeropad3D_CP_2152_elements(1115);
    -- CP-element group 7:  merge  fork  transition  place  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	1171 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	1126 
    -- CP-element group 7: 	1127 
    -- CP-element group 7: 	1129 
    -- CP-element group 7: 	1130 
    -- CP-element group 7: 	1132 
    -- CP-element group 7: 	1133 
    -- CP-element group 7:  members (27) 
      -- CP-element group 7: 	 branch_block_stmt_714/merge_stmt_4689__exit__
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/type_cast_4302/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/type_cast_4302/SplitProtocol/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/type_cast_4302/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/type_cast_4302/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/type_cast_4302/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/type_cast_4302/SplitProtocol/Update/cr
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4308/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4308/SplitProtocol/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4308/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4308/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4308/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4308/SplitProtocol/Update/cr
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/type_cast_4315/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/type_cast_4315/SplitProtocol/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/type_cast_4315/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/type_cast_4315/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/type_cast_4315/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/type_cast_4315/SplitProtocol/Update/cr
      -- 
    rr_13525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(7), ack => type_cast_4302_inst_req_0); -- 
    cr_13530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(7), ack => type_cast_4302_inst_req_1); -- 
    rr_13548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(7), ack => type_cast_4308_inst_req_0); -- 
    cr_13553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(7), ack => type_cast_4308_inst_req_1); -- 
    rr_13571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(7), ack => type_cast_4315_inst_req_0); -- 
    cr_13576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(7), ack => type_cast_4315_inst_req_1); -- 
    zeropad3D_CP_2152_elements(7) <= zeropad3D_CP_2152_elements(1171);
    -- CP-element group 8:  merge  fork  transition  place  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1233 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	1186 
    -- CP-element group 8: 	1187 
    -- CP-element group 8: 	1189 
    -- CP-element group 8: 	1190 
    -- CP-element group 8: 	1192 
    -- CP-element group 8: 	1193 
    -- CP-element group 8:  members (27) 
      -- CP-element group 8: 	 branch_block_stmt_714/merge_stmt_5246__exit__
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4879/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4879/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4879/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4879/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4879/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4879/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4883/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4883/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4883/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4883/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4883/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4883/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/type_cast_4873/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/type_cast_4873/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/type_cast_4873/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/type_cast_4873/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/type_cast_4873/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/type_cast_4873/SplitProtocol/Update/cr
      -- 
    rr_13961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(8), ack => type_cast_4879_inst_req_0); -- 
    cr_13966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(8), ack => type_cast_4879_inst_req_1); -- 
    rr_13984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(8), ack => type_cast_4883_inst_req_0); -- 
    cr_13989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(8), ack => type_cast_4883_inst_req_1); -- 
    rr_14007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(8), ack => type_cast_4873_inst_req_0); -- 
    cr_14012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(8), ack => type_cast_4873_inst_req_1); -- 
    zeropad3D_CP_2152_elements(8) <= zeropad3D_CP_2152_elements(1233);
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Sample/cra
      -- 
    cra_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_716_call_ack_0, ack => zeropad3D_CP_2152_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	35 
    -- CP-element group 10: 	36 
    -- CP-element group 10: 	37 
    -- CP-element group 10: 	38 
    -- CP-element group 10: 	39 
    -- CP-element group 10: 	40 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Update/cca
      -- 
    cca_2614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_716_call_ack_1, ack => zeropad3D_CP_2152_elements(10)); -- 
    -- CP-element group 11:  join  transition  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: 	37 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/word_access_start/$entry
      -- CP-element group 11: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/word_access_start/word_0/$entry
      -- CP-element group 11: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/word_access_start/word_0/rr
      -- 
    rr_2647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(11), ack => ptr_deref_727_load_0_req_0); -- 
    zeropad3D_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(0) & zeropad3D_CP_2152_elements(37);
      gj_zeropad3D_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/word_access_start/$exit
      -- CP-element group 12: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/word_access_start/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/word_access_start/word_0/ra
      -- 
    ra_2648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_727_load_0_ack_0, ack => zeropad3D_CP_2152_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (12) 
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/word_access_complete/$exit
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/word_access_complete/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/word_access_complete/word_0/ca
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/ptr_deref_727_Merge/$entry
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/ptr_deref_727_Merge/$exit
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/ptr_deref_727_Merge/merge_req
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/ptr_deref_727_Merge/merge_ack
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Sample/rr
      -- 
    ca_2659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_727_load_0_ack_1, ack => zeropad3D_CP_2152_elements(13)); -- 
    rr_2672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(13), ack => type_cast_731_inst_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Sample/ra
      -- 
    ra_2673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_0, ack => zeropad3D_CP_2152_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Update/ca
      -- 
    ca_2678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_1, ack => zeropad3D_CP_2152_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: 	15 
    -- CP-element group 16: 	40 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/STORE_row_high_733_Split/$entry
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/STORE_row_high_733_Split/$exit
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/STORE_row_high_733_Split/split_req
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/STORE_row_high_733_Split/split_ack
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/word_access_start/$entry
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/word_access_start/word_0/$entry
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/word_access_start/word_0/rr
      -- 
    rr_2699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(16), ack => STORE_row_high_733_store_0_req_0); -- 
    zeropad3D_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(0) & zeropad3D_CP_2152_elements(15) & zeropad3D_CP_2152_elements(40);
      gj_zeropad3D_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/word_access_start/word_0/ra
      -- 
    ra_2700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_row_high_733_store_0_ack_0, ack => zeropad3D_CP_2152_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	0 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	41 
    -- CP-element group 18:  members (5) 
      -- CP-element group 18: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/word_access_complete/word_0/ca
      -- 
    ca_2711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_row_high_733_store_0_ack_1, ack => zeropad3D_CP_2152_elements(18)); -- 
    -- CP-element group 19:  join  transition  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	0 
    -- CP-element group 19: 	38 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/word_access_start/$entry
      -- CP-element group 19: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/word_access_start/word_0/$entry
      -- CP-element group 19: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/word_access_start/word_0/rr
      -- 
    rr_2744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(19), ack => ptr_deref_746_load_0_req_0); -- 
    zeropad3D_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(0) & zeropad3D_CP_2152_elements(38);
      gj_zeropad3D_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/word_access_start/$exit
      -- CP-element group 20: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/word_access_start/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/word_access_start/word_0/ra
      -- 
    ra_2745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_746_load_0_ack_0, ack => zeropad3D_CP_2152_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (12) 
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/word_access_complete/$exit
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/word_access_complete/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/word_access_complete/word_0/ca
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/ptr_deref_746_Merge/$entry
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/ptr_deref_746_Merge/$exit
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/ptr_deref_746_Merge/merge_req
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/ptr_deref_746_Merge/merge_ack
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Sample/rr
      -- 
    ca_2756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_746_load_0_ack_1, ack => zeropad3D_CP_2152_elements(21)); -- 
    rr_2769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(21), ack => type_cast_750_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Sample/ra
      -- 
    ra_2770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_0, ack => zeropad3D_CP_2152_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Update/ca
      -- 
    ca_2775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_1, ack => zeropad3D_CP_2152_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: 	23 
    -- CP-element group 24: 	35 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/STORE_col_high_752_Split/$entry
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/STORE_col_high_752_Split/$exit
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/STORE_col_high_752_Split/split_req
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/STORE_col_high_752_Split/split_ack
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/word_access_start/$entry
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/word_access_start/word_0/$entry
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/word_access_start/word_0/rr
      -- 
    rr_2796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(24), ack => STORE_col_high_752_store_0_req_0); -- 
    zeropad3D_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(0) & zeropad3D_CP_2152_elements(23) & zeropad3D_CP_2152_elements(35);
      gj_zeropad3D_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/word_access_start/word_0/ra
      -- 
    ra_2797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_col_high_752_store_0_ack_0, ack => zeropad3D_CP_2152_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	0 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	41 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/word_access_complete/word_0/ca
      -- 
    ca_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_col_high_752_store_0_ack_1, ack => zeropad3D_CP_2152_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: 	39 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/word_access_start/$entry
      -- CP-element group 27: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/word_access_start/word_0/$entry
      -- CP-element group 27: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/word_access_start/word_0/rr
      -- 
    rr_2841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(27), ack => ptr_deref_765_load_0_req_0); -- 
    zeropad3D_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(0) & zeropad3D_CP_2152_elements(39);
      gj_zeropad3D_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (5) 
      -- CP-element group 28: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/word_access_start/$exit
      -- CP-element group 28: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/word_access_start/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/word_access_start/word_0/ra
      -- 
    ra_2842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_765_load_0_ack_0, ack => zeropad3D_CP_2152_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (12) 
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/word_access_complete/$exit
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/word_access_complete/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/word_access_complete/word_0/ca
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/ptr_deref_765_Merge/$entry
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/ptr_deref_765_Merge/$exit
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/ptr_deref_765_Merge/merge_req
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/ptr_deref_765_Merge/merge_ack
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Sample/rr
      -- 
    ca_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_765_load_0_ack_1, ack => zeropad3D_CP_2152_elements(29)); -- 
    rr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(29), ack => type_cast_769_inst_req_0); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Sample/ra
      -- 
    ra_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_769_inst_ack_0, ack => zeropad3D_CP_2152_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	0 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Update/ca
      -- 
    ca_2872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_769_inst_ack_1, ack => zeropad3D_CP_2152_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: 	31 
    -- CP-element group 32: 	36 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (9) 
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/STORE_depth_high_771_Split/$entry
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/STORE_depth_high_771_Split/$exit
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/STORE_depth_high_771_Split/split_req
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/STORE_depth_high_771_Split/split_ack
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/word_access_start/$entry
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/word_access_start/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/word_access_start/word_0/rr
      -- 
    rr_2893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(32), ack => STORE_depth_high_771_store_0_req_0); -- 
    zeropad3D_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(0) & zeropad3D_CP_2152_elements(31) & zeropad3D_CP_2152_elements(36);
      gj_zeropad3D_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/word_access_start/word_0/ra
      -- 
    ra_2894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_depth_high_771_store_0_ack_0, ack => zeropad3D_CP_2152_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	0 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	41 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/word_access_complete/word_0/ca
      -- 
    ca_2905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_depth_high_771_store_0_ack_1, ack => zeropad3D_CP_2152_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	10 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	24 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_STORE_col_high_752_delay
      -- 
    -- Element group zeropad3D_CP_2152_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(10), ack => zeropad3D_CP_2152_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  transition  delay-element  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	10 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	32 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_STORE_depth_high_771_delay
      -- 
    -- Element group zeropad3D_CP_2152_elements(36) is a control-delay.
    cp_element_36_delay: control_delay_element  generic map(name => " 36_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(10), ack => zeropad3D_CP_2152_elements(36), clk => clk, reset =>reset);
    -- CP-element group 37:  transition  delay-element  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	10 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	11 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_ptr_deref_727_delay
      -- 
    -- Element group zeropad3D_CP_2152_elements(37) is a control-delay.
    cp_element_37_delay: control_delay_element  generic map(name => " 37_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(10), ack => zeropad3D_CP_2152_elements(37), clk => clk, reset =>reset);
    -- CP-element group 38:  transition  delay-element  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	10 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	19 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_ptr_deref_746_delay
      -- 
    -- Element group zeropad3D_CP_2152_elements(38) is a control-delay.
    cp_element_38_delay: control_delay_element  generic map(name => " 38_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(10), ack => zeropad3D_CP_2152_elements(38), clk => clk, reset =>reset);
    -- CP-element group 39:  transition  delay-element  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	10 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	27 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_ptr_deref_765_delay
      -- 
    -- Element group zeropad3D_CP_2152_elements(39) is a control-delay.
    cp_element_39_delay: control_delay_element  generic map(name => " 39_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(10), ack => zeropad3D_CP_2152_elements(39), clk => clk, reset =>reset);
    -- CP-element group 40:  transition  delay-element  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	10 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	16 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_STORE_row_high_733_delay
      -- 
    -- Element group zeropad3D_CP_2152_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(10), ack => zeropad3D_CP_2152_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  fork  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: 	26 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: 	43 
    -- CP-element group 41: 	44 
    -- CP-element group 41: 	45 
    -- CP-element group 41: 	46 
    -- CP-element group 41: 	47 
    -- CP-element group 41: 	48 
    -- CP-element group 41: 	49 
    -- CP-element group 41: 	50 
    -- CP-element group 41: 	51 
    -- CP-element group 41: 	53 
    -- CP-element group 41: 	55 
    -- CP-element group 41: 	57 
    -- CP-element group 41:  members (101) 
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896__entry__
      -- CP-element group 41: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773__exit__
      -- CP-element group 41: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/word_access_start/word_0/rr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/word_access_start/word_0/rr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/word_access_start/word_0/rr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_address_resized
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_addr_resize/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_addr_resize/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_addr_resize/base_resize_req
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_addr_resize/base_resize_ack
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_word_addrgen/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_word_addrgen/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_word_addrgen/root_register_req
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_word_addrgen/root_register_ack
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/word_access_start/word_0/rr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_address_resized
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_addr_resize/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_addr_resize/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_addr_resize/base_resize_req
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_addr_resize/base_resize_ack
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_word_addrgen/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_word_addrgen/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_word_addrgen/root_register_req
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_word_addrgen/root_register_ack
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/word_access_start/word_0/rr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Update/cr
      -- 
    rr_2930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => LOAD_pad_776_load_0_req_0); -- 
    cr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => LOAD_pad_776_load_0_req_1); -- 
    rr_2963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => LOAD_depth_high_779_load_0_req_0); -- 
    cr_2974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => LOAD_depth_high_779_load_0_req_1); -- 
    rr_2996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => LOAD_col_high_782_load_0_req_0); -- 
    cr_3007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => LOAD_col_high_782_load_0_req_1); -- 
    rr_3046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => ptr_deref_794_load_0_req_0); -- 
    cr_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => ptr_deref_794_load_0_req_1); -- 
    rr_3096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => ptr_deref_806_load_0_req_0); -- 
    cr_3107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => ptr_deref_806_load_0_req_1); -- 
    cr_3126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => type_cast_810_inst_req_1); -- 
    cr_3140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => type_cast_814_inst_req_1); -- 
    cr_3154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => type_cast_854_inst_req_1); -- 
    zeropad3D_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(18) & zeropad3D_CP_2152_elements(26) & zeropad3D_CP_2152_elements(34);
      gj_zeropad3D_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/word_access_start/$exit
      -- CP-element group 42: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/word_access_start/word_0/ra
      -- 
    ra_2931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_776_load_0_ack_0, ack => zeropad3D_CP_2152_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	56 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/word_access_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/word_access_complete/word_0/ca
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/LOAD_pad_776_Merge/$entry
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/LOAD_pad_776_Merge/$exit
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/LOAD_pad_776_Merge/merge_req
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/LOAD_pad_776_Merge/merge_ack
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Sample/rr
      -- 
    ca_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_776_load_0_ack_1, ack => zeropad3D_CP_2152_elements(43)); -- 
    rr_3149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(43), ack => type_cast_854_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	41 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/word_access_start/$exit
      -- CP-element group 44: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/word_access_start/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/word_access_start/word_0/ra
      -- 
    ra_2964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_779_load_0_ack_0, ack => zeropad3D_CP_2152_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	41 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	52 
    -- CP-element group 45:  members (12) 
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/word_access_complete/$exit
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/word_access_complete/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/word_access_complete/word_0/ca
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/LOAD_depth_high_779_Merge/$entry
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/LOAD_depth_high_779_Merge/$exit
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/LOAD_depth_high_779_Merge/merge_req
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/LOAD_depth_high_779_Merge/merge_ack
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Sample/rr
      -- 
    ca_2975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_779_load_0_ack_1, ack => zeropad3D_CP_2152_elements(45)); -- 
    rr_3121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(45), ack => type_cast_810_inst_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	41 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/word_access_start/$exit
      -- CP-element group 46: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/word_access_start/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/word_access_start/word_0/ra
      -- 
    ra_2997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_782_load_0_ack_0, ack => zeropad3D_CP_2152_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	41 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	54 
    -- CP-element group 47:  members (12) 
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/word_access_complete/$exit
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/word_access_complete/word_0/$exit
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/word_access_complete/word_0/ca
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/LOAD_col_high_782_Merge/$entry
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/LOAD_col_high_782_Merge/$exit
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/LOAD_col_high_782_Merge/merge_req
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/LOAD_col_high_782_Merge/merge_ack
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Sample/rr
      -- 
    ca_3008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_782_load_0_ack_1, ack => zeropad3D_CP_2152_elements(47)); -- 
    rr_3135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(47), ack => type_cast_814_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	41 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/word_access_start/$exit
      -- CP-element group 48: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/word_access_start/word_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/word_access_start/word_0/ra
      -- 
    ra_3047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_794_load_0_ack_0, ack => zeropad3D_CP_2152_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	41 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (9) 
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/word_access_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/word_access_complete/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/word_access_complete/word_0/ca
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/ptr_deref_794_Merge/$entry
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/ptr_deref_794_Merge/$exit
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/ptr_deref_794_Merge/merge_req
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/ptr_deref_794_Merge/merge_ack
      -- 
    ca_3058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_794_load_0_ack_1, ack => zeropad3D_CP_2152_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/word_access_start/$exit
      -- CP-element group 50: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/word_access_start/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/word_access_start/word_0/ra
      -- 
    ra_3097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_806_load_0_ack_0, ack => zeropad3D_CP_2152_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	41 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	58 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/word_access_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/word_access_complete/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/word_access_complete/word_0/ca
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/ptr_deref_806_Merge/$entry
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/ptr_deref_806_Merge/$exit
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/ptr_deref_806_Merge/merge_req
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/ptr_deref_806_Merge/merge_ack
      -- 
    ca_3108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_806_load_0_ack_1, ack => zeropad3D_CP_2152_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	45 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Sample/ra
      -- 
    ra_3122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_810_inst_ack_0, ack => zeropad3D_CP_2152_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	41 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	58 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Update/ca
      -- 
    ca_3127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_810_inst_ack_1, ack => zeropad3D_CP_2152_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	47 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Sample/ra
      -- 
    ra_3136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_814_inst_ack_0, ack => zeropad3D_CP_2152_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	41 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Update/ca
      -- 
    ca_3141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_814_inst_ack_1, ack => zeropad3D_CP_2152_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Sample/ra
      -- 
    ra_3150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_0, ack => zeropad3D_CP_2152_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	41 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Update/ca
      -- 
    ca_3155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_1, ack => zeropad3D_CP_2152_elements(57)); -- 
    -- CP-element group 58:  join  fork  transition  place  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	49 
    -- CP-element group 58: 	51 
    -- CP-element group 58: 	53 
    -- CP-element group 58: 	55 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	780 
    -- CP-element group 58: 	781 
    -- CP-element group 58: 	782 
    -- CP-element group 58:  members (10) 
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody
      -- CP-element group 58: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896__exit__
      -- CP-element group 58: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/$exit
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/$entry
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_913/$entry
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/$entry
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_906/$entry
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/$entry
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_899/$entry
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(49) & zeropad3D_CP_2152_elements(51) & zeropad3D_CP_2152_elements(53) & zeropad3D_CP_2152_elements(55) & zeropad3D_CP_2152_elements(57);
      gj_zeropad3D_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	798 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Sample/ra
      -- 
    ra_3167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_924_inst_ack_0, ack => zeropad3D_CP_2152_elements(59)); -- 
    -- CP-element group 60:  branch  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	798 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (13) 
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933__entry__
      -- CP-element group 60: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932__exit__
      -- CP-element group 60: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/$exit
      -- CP-element group 60: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933_dead_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933_eval_test/$entry
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933_eval_test/$exit
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933_eval_test/branch_req
      -- CP-element group 60: 	 branch_block_stmt_714/R_cmp_934_place
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933_if_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933_else_link/$entry
      -- 
    ca_3172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_924_inst_ack_1, ack => zeropad3D_CP_2152_elements(60)); -- 
    branch_req_3180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(60), ack => if_stmt_933_branch_req_0); -- 
    -- CP-element group 61:  transition  place  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	799 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 branch_block_stmt_714/whilex_xbody_ifx_xthen
      -- CP-element group 61: 	 branch_block_stmt_714/if_stmt_933_if_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_714/if_stmt_933_if_link/if_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_714/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 61: 	 branch_block_stmt_714/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- 
    if_choice_transition_3185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_933_branch_ack_1, ack => zeropad3D_CP_2152_elements(61)); -- 
    -- CP-element group 62:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62: 	66 
    -- CP-element group 62:  members (27) 
      -- CP-element group 62: 	 branch_block_stmt_714/merge_stmt_939__exit__
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964__entry__
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/word_access_start/word_0/rr
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/word_access_complete/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_update_start_
      -- CP-element group 62: 	 branch_block_stmt_714/whilex_xbody_lorx_xlhsx_xfalse
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_update_start_
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/word_access_start/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/word_access_complete/word_0/cr
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/word_access_start/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/if_stmt_933_else_link/else_choice_transition
      -- CP-element group 62: 	 branch_block_stmt_714/if_stmt_933_else_link/$exit
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/word_access_complete/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/merge_stmt_939_PhiReqMerge
      -- CP-element group 62: 	 branch_block_stmt_714/merge_stmt_939_PhiAck/dummy
      -- CP-element group 62: 	 branch_block_stmt_714/merge_stmt_939_PhiAck/$exit
      -- CP-element group 62: 	 branch_block_stmt_714/merge_stmt_939_PhiAck/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_714/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$entry
      -- 
    else_choice_transition_3189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_933_branch_ack_0, ack => zeropad3D_CP_2152_elements(62)); -- 
    rr_3210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(62), ack => LOAD_row_high_941_load_0_req_0); -- 
    cr_3221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(62), ack => LOAD_row_high_941_load_0_req_1); -- 
    cr_3240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(62), ack => type_cast_945_inst_req_1); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/word_access_start/word_0/ra
      -- CP-element group 63: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/word_access_start/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/word_access_start/$exit
      -- CP-element group 63: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/$exit
      -- 
    ra_3211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_941_load_0_ack_0, ack => zeropad3D_CP_2152_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (12) 
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/LOAD_row_high_941_Merge/merge_req
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/word_access_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/LOAD_row_high_941_Merge/merge_ack
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/LOAD_row_high_941_Merge/$exit
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/LOAD_row_high_941_Merge/$entry
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/word_access_complete/word_0/ca
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/word_access_complete/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Sample/$entry
      -- 
    ca_3222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_941_load_0_ack_1, ack => zeropad3D_CP_2152_elements(64)); -- 
    rr_3235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(64), ack => type_cast_945_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Sample/ra
      -- CP-element group 65: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Sample/$exit
      -- 
    ra_3236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_945_inst_ack_0, ack => zeropad3D_CP_2152_elements(65)); -- 
    -- CP-element group 66:  branch  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	62 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (13) 
      -- CP-element group 66: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964__exit__
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965__entry__
      -- CP-element group 66: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_714/R_cmp56_966_place
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965_else_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/$exit
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Update/$exit
      -- 
    ca_3241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_945_inst_ack_1, ack => zeropad3D_CP_2152_elements(66)); -- 
    branch_req_3249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(66), ack => if_stmt_965_branch_req_0); -- 
    -- CP-element group 67:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: 	70 
    -- CP-element group 67:  members (18) 
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_714/merge_stmt_971__exit__
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983__entry__
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_714/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse58
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_update_start_
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/$entry
      -- CP-element group 67: 	 branch_block_stmt_714/if_stmt_965_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_714/if_stmt_965_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_714/merge_stmt_971_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_714/merge_stmt_971_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_714/merge_stmt_971_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_714/merge_stmt_971_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_714/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse58_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_714/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse58_PhiReq/$entry
      -- 
    if_choice_transition_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_965_branch_ack_1, ack => zeropad3D_CP_2152_elements(67)); -- 
    cr_3276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(67), ack => type_cast_975_inst_req_1); -- 
    rr_3271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(67), ack => type_cast_975_inst_req_0); -- 
    -- CP-element group 68:  transition  place  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	799 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 branch_block_stmt_714/lorx_xlhsx_xfalse_ifx_xthen
      -- CP-element group 68: 	 branch_block_stmt_714/if_stmt_965_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_714/if_stmt_965_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_714/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_714/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_3258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_965_branch_ack_0, ack => zeropad3D_CP_2152_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_sample_completed_
      -- 
    ra_3272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_975_inst_ack_0, ack => zeropad3D_CP_2152_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	67 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983__exit__
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984__entry__
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/$exit
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984_else_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_714/R_cmp63_985_place
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984_eval_test/$entry
      -- 
    ca_3277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_975_inst_ack_1, ack => zeropad3D_CP_2152_elements(70)); -- 
    branch_req_3285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(70), ack => if_stmt_984_branch_req_0); -- 
    -- CP-element group 71:  transition  place  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	799 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_714/lorx_xlhsx_xfalse58_ifx_xthen
      -- CP-element group 71: 	 branch_block_stmt_714/if_stmt_984_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_714/if_stmt_984_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_714/lorx_xlhsx_xfalse58_ifx_xthen_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_714/lorx_xlhsx_xfalse58_ifx_xthen_PhiReq/$entry
      -- 
    if_choice_transition_3290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_984_branch_ack_1, ack => zeropad3D_CP_2152_elements(71)); -- 
    -- CP-element group 72:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: 	74 
    -- CP-element group 72: 	76 
    -- CP-element group 72:  members (27) 
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015__entry__
      -- CP-element group 72: 	 branch_block_stmt_714/merge_stmt_990__exit__
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Update/cr
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_update_start_
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/word_access_complete/word_0/cr
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/word_access_complete/word_0/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/word_access_complete/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/word_access_start/word_0/rr
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/word_access_start/word_0/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/word_access_start/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_root_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_word_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_update_start_
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/lorx_xlhsx_xfalse58_lorx_xlhsx_xfalse65
      -- CP-element group 72: 	 branch_block_stmt_714/if_stmt_984_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_714/if_stmt_984_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_714/merge_stmt_990_PhiAck/dummy
      -- CP-element group 72: 	 branch_block_stmt_714/merge_stmt_990_PhiAck/$exit
      -- CP-element group 72: 	 branch_block_stmt_714/merge_stmt_990_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/merge_stmt_990_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_714/lorx_xlhsx_xfalse58_lorx_xlhsx_xfalse65_PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_714/lorx_xlhsx_xfalse58_lorx_xlhsx_xfalse65_PhiReq/$entry
      -- 
    else_choice_transition_3294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_984_branch_ack_0, ack => zeropad3D_CP_2152_elements(72)); -- 
    cr_3345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(72), ack => type_cast_996_inst_req_1); -- 
    cr_3326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(72), ack => LOAD_col_high_992_load_0_req_1); -- 
    rr_3315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(72), ack => LOAD_col_high_992_load_0_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/word_access_start/word_0/ra
      -- CP-element group 73: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/word_access_start/word_0/$exit
      -- CP-element group 73: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/word_access_start/$exit
      -- CP-element group 73: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_sample_completed_
      -- 
    ra_3316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_992_load_0_ack_0, ack => zeropad3D_CP_2152_elements(73)); -- 
    -- CP-element group 74:  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (12) 
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/LOAD_col_high_992_Merge/merge_ack
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/LOAD_col_high_992_Merge/merge_req
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/LOAD_col_high_992_Merge/$exit
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/LOAD_col_high_992_Merge/$entry
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/word_access_complete/word_0/ca
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/word_access_complete/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/word_access_complete/$exit
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_update_completed_
      -- 
    ca_3327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_992_load_0_ack_1, ack => zeropad3D_CP_2152_elements(74)); -- 
    rr_3340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(74), ack => type_cast_996_inst_req_0); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_sample_completed_
      -- 
    ra_3341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_996_inst_ack_0, ack => zeropad3D_CP_2152_elements(75)); -- 
    -- CP-element group 76:  branch  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	72 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (13) 
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016__entry__
      -- CP-element group 76: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015__exit__
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016_else_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016_if_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_714/R_cmp74_1017_place
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016_eval_test/branch_req
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016_eval_test/$exit
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016_eval_test/$entry
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016_dead_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/$exit
      -- 
    ca_3346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_996_inst_ack_1, ack => zeropad3D_CP_2152_elements(76)); -- 
    branch_req_3354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(76), ack => if_stmt_1016_branch_req_0); -- 
    -- CP-element group 77:  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	93 
    -- CP-element group 77: 	94 
    -- CP-element group 77: 	96 
    -- CP-element group 77: 	98 
    -- CP-element group 77: 	100 
    -- CP-element group 77: 	102 
    -- CP-element group 77: 	104 
    -- CP-element group 77: 	106 
    -- CP-element group 77: 	108 
    -- CP-element group 77: 	111 
    -- CP-element group 77:  members (46) 
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186__entry__
      -- CP-element group 77: 	 branch_block_stmt_714/merge_stmt_1081__exit__
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/if_stmt_1016_if_link/$exit
      -- CP-element group 77: 	 branch_block_stmt_714/if_stmt_1016_if_link/if_choice_transition
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/lorx_xlhsx_xfalse65_ifx_xelse
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Update/req
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_complete/req
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_update_start
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_update_start
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Update/req
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_complete/req
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_714/merge_stmt_1081_PhiAck/dummy
      -- CP-element group 77: 	 branch_block_stmt_714/merge_stmt_1081_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_714/merge_stmt_1081_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/merge_stmt_1081_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_714/lorx_xlhsx_xfalse65_ifx_xelse_PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_714/lorx_xlhsx_xfalse65_ifx_xelse_PhiReq/$entry
      -- 
    if_choice_transition_3359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1016_branch_ack_1, ack => zeropad3D_CP_2152_elements(77)); -- 
    cr_3522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => type_cast_1085_inst_req_1); -- 
    rr_3517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => type_cast_1085_inst_req_0); -- 
    cr_3627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => ptr_deref_1160_load_0_req_1); -- 
    req_3567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => array_obj_ref_1155_index_offset_req_1); -- 
    cr_3536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => type_cast_1149_inst_req_1); -- 
    req_3582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => addr_of_1156_final_reg_req_1); -- 
    cr_3646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => type_cast_1174_inst_req_1); -- 
    req_3677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => array_obj_ref_1180_index_offset_req_1); -- 
    req_3692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => addr_of_1181_final_reg_req_1); -- 
    cr_3742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => ptr_deref_1184_store_0_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	799 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_714/if_stmt_1016_else_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_714/if_stmt_1016_else_link/else_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_714/lorx_xlhsx_xfalse65_ifx_xthen
      -- CP-element group 78: 	 branch_block_stmt_714/lorx_xlhsx_xfalse65_ifx_xthen_PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_714/lorx_xlhsx_xfalse65_ifx_xthen_PhiReq/$entry
      -- 
    else_choice_transition_3363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1016_branch_ack_0, ack => zeropad3D_CP_2152_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	799 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Sample/ra
      -- CP-element group 79: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_sample_completed_
      -- 
    ra_3377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1026_inst_ack_0, ack => zeropad3D_CP_2152_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	799 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_update_completed_
      -- 
    ca_3382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1026_inst_ack_1, ack => zeropad3D_CP_2152_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	799 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Sample/$exit
      -- 
    ra_3391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1031_inst_ack_0, ack => zeropad3D_CP_2152_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	799 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_update_completed_
      -- 
    ca_3396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1031_inst_ack_1, ack => zeropad3D_CP_2152_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_sample_start_
      -- 
    rr_3404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(83), ack => type_cast_1066_inst_req_0); -- 
    zeropad3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(80) & zeropad3D_CP_2152_elements(82);
      gj_zeropad3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_sample_completed_
      -- 
    ra_3405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1066_inst_ack_0, ack => zeropad3D_CP_2152_elements(84)); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	799 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (16) 
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_resize_1/$exit
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_resize_1/index_resize_req
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_resize_1/index_resize_ack
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_resize_1/$entry
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_computed_1
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_scaled_1
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_resized_1
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Update/ca
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Sample/req
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_scale_1/scale_rename_ack
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_scale_1/scale_rename_req
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_scale_1/$exit
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_scale_1/$entry
      -- 
    ca_3410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1066_inst_ack_1, ack => zeropad3D_CP_2152_elements(85)); -- 
    req_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(85), ack => array_obj_ref_1072_index_offset_req_0); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	92 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Sample/ack
      -- CP-element group 86: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_sample_complete
      -- 
    ack_3436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1072_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(86)); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	799 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (11) 
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_offset_calculated
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_root_address_calculated
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_request/req
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_request/$entry
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_base_plus_offset/sum_rename_ack
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_base_plus_offset/sum_rename_req
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_base_plus_offset/$exit
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_base_plus_offset/$entry
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Update/ack
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Update/$exit
      -- 
    ack_3441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1072_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(87)); -- 
    req_3450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(87), ack => addr_of_1073_final_reg_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_request/ack
      -- CP-element group 88: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_request/$exit
      -- 
    ack_3451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1073_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(88)); -- 
    -- CP-element group 89:  join  fork  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	799 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (28) 
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_word_addrgen/root_register_ack
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/word_access_start/$entry
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_plus_offset/sum_rename_ack
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_word_addrgen/$entry
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/word_access_start/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_word_addrgen/$exit
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_plus_offset/sum_rename_req
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_plus_offset/$exit
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_plus_offset/$entry
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_addr_resize/base_resize_ack
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_addr_resize/base_resize_req
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_addr_resize/$exit
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_addr_resize/$entry
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_address_resized
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_root_address_calculated
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/ptr_deref_1076_Split/split_ack
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_word_address_calculated
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_address_calculated
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_complete/ack
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/ptr_deref_1076_Split/split_req
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_complete/$exit
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/ptr_deref_1076_Split/$exit
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_word_addrgen/root_register_req
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/ptr_deref_1076_Split/$entry
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/word_access_start/word_0/rr
      -- 
    ack_3456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1073_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(89)); -- 
    rr_3494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(89), ack => ptr_deref_1076_store_0_req_0); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/word_access_start/$exit
      -- CP-element group 90: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/word_access_start/word_0/$exit
      -- CP-element group 90: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/word_access_start/word_0/ra
      -- 
    ra_3495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1076_store_0_ack_0, ack => zeropad3D_CP_2152_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	799 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/word_access_complete/word_0/ca
      -- CP-element group 91: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/word_access_complete/word_0/$exit
      -- CP-element group 91: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/word_access_complete/$exit
      -- CP-element group 91: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/$exit
      -- 
    ca_3506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1076_store_0_ack_1, ack => zeropad3D_CP_2152_elements(91)); -- 
    -- CP-element group 92:  join  transition  place  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	86 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	800 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079__exit__
      -- CP-element group 92: 	 branch_block_stmt_714/ifx_xthen_ifx_xend
      -- CP-element group 92: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/$exit
      -- CP-element group 92: 	 branch_block_stmt_714/ifx_xthen_ifx_xend_PhiReq/$exit
      -- CP-element group 92: 	 branch_block_stmt_714/ifx_xthen_ifx_xend_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(86) & zeropad3D_CP_2152_elements(91);
      gj_zeropad3D_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	77 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_sample_completed_
      -- 
    ra_3518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1085_inst_ack_0, ack => zeropad3D_CP_2152_elements(93)); -- 
    -- CP-element group 94:  fork  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	77 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94: 	103 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Update/ca
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Sample/rr
      -- 
    ca_3523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1085_inst_ack_1, ack => zeropad3D_CP_2152_elements(94)); -- 
    rr_3531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(94), ack => type_cast_1149_inst_req_0); -- 
    rr_3641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(94), ack => type_cast_1174_inst_req_0); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Sample/$exit
      -- 
    ra_3532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1149_inst_ack_0, ack => zeropad3D_CP_2152_elements(95)); -- 
    -- CP-element group 96:  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	77 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (16) 
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_computed_1
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_resize_1/$entry
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_resize_1/$exit
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_scaled_1
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_resized_1
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Sample/req
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_scale_1/scale_rename_ack
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_scale_1/scale_rename_req
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_scale_1/$exit
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_scale_1/$entry
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_resize_1/index_resize_ack
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_resize_1/index_resize_req
      -- 
    ca_3537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1149_inst_ack_1, ack => zeropad3D_CP_2152_elements(96)); -- 
    req_3562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(96), ack => array_obj_ref_1155_index_offset_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	112 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Sample/ack
      -- CP-element group 97: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_sample_complete
      -- 
    ack_3563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1155_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	77 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (11) 
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_request/req
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_request/$entry
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_base_plus_offset/sum_rename_ack
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_base_plus_offset/sum_rename_req
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_offset_calculated
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_root_address_calculated
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_base_plus_offset/$exit
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_base_plus_offset/$entry
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Update/ack
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_sample_start_
      -- 
    ack_3568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1155_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(98)); -- 
    req_3577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(98), ack => addr_of_1156_final_reg_req_0); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_request/ack
      -- CP-element group 99: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_request/$exit
      -- CP-element group 99: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_sample_completed_
      -- 
    ack_3578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1156_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	77 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (24) 
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_plus_offset/sum_rename_req
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_plus_offset/$exit
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_plus_offset/$entry
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/word_access_start/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_addr_resize/base_resize_ack
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_addr_resize/base_resize_req
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_word_addrgen/$exit
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_addr_resize/$exit
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_addr_resize/$entry
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_address_resized
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_root_address_calculated
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_word_address_calculated
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_address_calculated
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_word_addrgen/$entry
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/word_access_start/word_0/rr
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/word_access_start/$entry
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_complete/ack
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_complete/$exit
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_word_addrgen/root_register_ack
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_word_addrgen/root_register_req
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_plus_offset/sum_rename_ack
      -- 
    ack_3583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1156_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(100)); -- 
    rr_3616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(100), ack => ptr_deref_1160_load_0_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/word_access_start/word_0/ra
      -- CP-element group 101: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/word_access_start/$exit
      -- CP-element group 101: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/word_access_start/word_0/$exit
      -- 
    ra_3617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1160_load_0_ack_0, ack => zeropad3D_CP_2152_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	77 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	109 
    -- CP-element group 102:  members (9) 
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/ptr_deref_1160_Merge/$exit
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/ptr_deref_1160_Merge/$entry
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/word_access_complete/word_0/ca
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/word_access_complete/word_0/$exit
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/ptr_deref_1160_Merge/merge_ack
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/word_access_complete/$exit
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/ptr_deref_1160_Merge/merge_req
      -- 
    ca_3628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1160_load_0_ack_1, ack => zeropad3D_CP_2152_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	94 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Sample/ra
      -- 
    ra_3642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1174_inst_ack_0, ack => zeropad3D_CP_2152_elements(103)); -- 
    -- CP-element group 104:  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	77 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (16) 
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_resized_1
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_scaled_1
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_computed_1
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_resize_1/$entry
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_resize_1/$exit
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_resize_1/index_resize_req
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_resize_1/index_resize_ack
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_scale_1/$entry
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_scale_1/$exit
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_scale_1/scale_rename_req
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_scale_1/scale_rename_ack
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Sample/req
      -- 
    ca_3647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1174_inst_ack_1, ack => zeropad3D_CP_2152_elements(104)); -- 
    req_3672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(104), ack => array_obj_ref_1180_index_offset_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	112 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_sample_complete
      -- CP-element group 105: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Sample/ack
      -- 
    ack_3673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1180_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	77 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (11) 
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_request/$entry
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_root_address_calculated
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_offset_calculated
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Update/ack
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_base_plus_offset/$entry
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_base_plus_offset/$exit
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_base_plus_offset/sum_rename_req
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_base_plus_offset/sum_rename_ack
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_request/req
      -- 
    ack_3678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1180_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(106)); -- 
    req_3687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(106), ack => addr_of_1181_final_reg_req_0); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_request/$exit
      -- CP-element group 107: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_request/ack
      -- 
    ack_3688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1181_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(107)); -- 
    -- CP-element group 108:  fork  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	77 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (19) 
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_complete/$exit
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_complete/ack
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_address_calculated
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_word_address_calculated
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_root_address_calculated
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_address_resized
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_addr_resize/$entry
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_addr_resize/$exit
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_addr_resize/base_resize_req
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_addr_resize/base_resize_ack
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_plus_offset/$entry
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_plus_offset/$exit
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_plus_offset/sum_rename_req
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_plus_offset/sum_rename_ack
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_word_addrgen/$entry
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_word_addrgen/$exit
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_word_addrgen/root_register_req
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_word_addrgen/root_register_ack
      -- 
    ack_3693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1181_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	102 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (9) 
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/ptr_deref_1184_Split/$entry
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/ptr_deref_1184_Split/$exit
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/ptr_deref_1184_Split/split_req
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/ptr_deref_1184_Split/split_ack
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/word_access_start/$entry
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/word_access_start/word_0/$entry
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/word_access_start/word_0/rr
      -- 
    rr_3731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(109), ack => ptr_deref_1184_store_0_req_0); -- 
    zeropad3D_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(102) & zeropad3D_CP_2152_elements(108);
      gj_zeropad3D_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/word_access_start/$exit
      -- CP-element group 110: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/word_access_start/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/word_access_start/word_0/ra
      -- 
    ra_3732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1184_store_0_ack_0, ack => zeropad3D_CP_2152_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	77 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/word_access_complete/$exit
      -- CP-element group 111: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/word_access_complete/word_0/$exit
      -- CP-element group 111: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/word_access_complete/word_0/ca
      -- 
    ca_3743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1184_store_0_ack_1, ack => zeropad3D_CP_2152_elements(111)); -- 
    -- CP-element group 112:  join  transition  place  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	97 
    -- CP-element group 112: 	105 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	800 
    -- CP-element group 112:  members (5) 
      -- CP-element group 112: 	 branch_block_stmt_714/ifx_xelse_ifx_xend
      -- CP-element group 112: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186__exit__
      -- CP-element group 112: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/$exit
      -- CP-element group 112: 	 branch_block_stmt_714/ifx_xelse_ifx_xend_PhiReq/$exit
      -- CP-element group 112: 	 branch_block_stmt_714/ifx_xelse_ifx_xend_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(97) & zeropad3D_CP_2152_elements(105) & zeropad3D_CP_2152_elements(111);
      gj_zeropad3D_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	800 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Sample/ra
      -- 
    ra_3755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1192_inst_ack_0, ack => zeropad3D_CP_2152_elements(113)); -- 
    -- CP-element group 114:  branch  transition  place  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	800 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (13) 
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207__entry__
      -- CP-element group 114: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206__exit__
      -- CP-element group 114: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/$exit
      -- CP-element group 114: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Update/ca
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207_dead_link/$entry
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207_eval_test/$entry
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207_eval_test/$exit
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207_eval_test/branch_req
      -- CP-element group 114: 	 branch_block_stmt_714/R_cmp143_1208_place
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207_if_link/$entry
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207_else_link/$entry
      -- 
    ca_3760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1192_inst_ack_1, ack => zeropad3D_CP_2152_elements(114)); -- 
    branch_req_3768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(114), ack => if_stmt_1207_branch_req_0); -- 
    -- CP-element group 115:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	809 
    -- CP-element group 115: 	810 
    -- CP-element group 115: 	812 
    -- CP-element group 115: 	813 
    -- CP-element group 115: 	815 
    -- CP-element group 115: 	816 
    -- CP-element group 115:  members (40) 
      -- CP-element group 115: 	 branch_block_stmt_714/assign_stmt_1219__entry__
      -- CP-element group 115: 	 branch_block_stmt_714/merge_stmt_1213__exit__
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184
      -- CP-element group 115: 	 branch_block_stmt_714/assign_stmt_1219__exit__
      -- CP-element group 115: 	 branch_block_stmt_714/if_stmt_1207_if_link/$exit
      -- CP-element group 115: 	 branch_block_stmt_714/if_stmt_1207_if_link/if_choice_transition
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xend_ifx_xthen145
      -- CP-element group 115: 	 branch_block_stmt_714/assign_stmt_1219/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/assign_stmt_1219/$exit
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Update/cr
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/merge_stmt_1213_PhiAck/dummy
      -- CP-element group 115: 	 branch_block_stmt_714/merge_stmt_1213_PhiAck/$exit
      -- CP-element group 115: 	 branch_block_stmt_714/merge_stmt_1213_PhiAck/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/merge_stmt_1213_PhiReqMerge
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Update/cr
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xend_ifx_xthen145_PhiReq/$exit
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xend_ifx_xthen145_PhiReq/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Update/cr
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Sample/rr
      -- 
    if_choice_transition_3773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1207_branch_ack_1, ack => zeropad3D_CP_2152_elements(115)); -- 
    rr_11276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(115), ack => type_cast_1325_inst_req_0); -- 
    cr_11304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(115), ack => type_cast_1312_inst_req_1); -- 
    rr_11299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(115), ack => type_cast_1312_inst_req_0); -- 
    cr_11258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(115), ack => type_cast_1316_inst_req_1); -- 
    cr_11281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(115), ack => type_cast_1325_inst_req_1); -- 
    rr_11253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(115), ack => type_cast_1316_inst_req_0); -- 
    -- CP-element group 116:  fork  transition  place  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	118 
    -- CP-element group 116: 	119 
    -- CP-element group 116: 	120 
    -- CP-element group 116: 	122 
    -- CP-element group 116: 	125 
    -- CP-element group 116: 	127 
    -- CP-element group 116: 	128 
    -- CP-element group 116: 	129 
    -- CP-element group 116: 	131 
    -- CP-element group 116:  members (54) 
      -- CP-element group 116: 	 branch_block_stmt_714/merge_stmt_1221__exit__
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299__entry__
      -- CP-element group 116: 	 branch_block_stmt_714/if_stmt_1207_else_link/$exit
      -- CP-element group 116: 	 branch_block_stmt_714/if_stmt_1207_else_link/else_choice_transition
      -- CP-element group 116: 	 branch_block_stmt_714/ifx_xend_ifx_xelse150
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_word_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_root_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/word_access_start/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/word_access_start/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/word_access_start/word_0/rr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/word_access_complete/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/word_access_complete/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/word_access_complete/word_0/cr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_word_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_root_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/word_access_start/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/word_access_start/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/word_access_start/word_0/rr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/word_access_complete/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/word_access_complete/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/word_access_complete/word_0/cr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_714/merge_stmt_1221_PhiAck/dummy
      -- CP-element group 116: 	 branch_block_stmt_714/merge_stmt_1221_PhiAck/$exit
      -- CP-element group 116: 	 branch_block_stmt_714/merge_stmt_1221_PhiAck/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/merge_stmt_1221_PhiReqMerge
      -- CP-element group 116: 	 branch_block_stmt_714/ifx_xend_ifx_xelse150_PhiReq/$exit
      -- CP-element group 116: 	 branch_block_stmt_714/ifx_xend_ifx_xelse150_PhiReq/$entry
      -- 
    else_choice_transition_3777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1207_branch_ack_0, ack => zeropad3D_CP_2152_elements(116)); -- 
    rr_3793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => type_cast_1231_inst_req_0); -- 
    cr_3798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => type_cast_1231_inst_req_1); -- 
    rr_3815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => LOAD_col_high_1234_load_0_req_0); -- 
    cr_3826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => LOAD_col_high_1234_load_0_req_1); -- 
    cr_3845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => type_cast_1238_inst_req_1); -- 
    cr_3859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => type_cast_1258_inst_req_1); -- 
    cr_3873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => type_cast_1275_inst_req_1); -- 
    rr_3890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => LOAD_row_high_1278_load_0_req_0); -- 
    cr_3901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => LOAD_row_high_1278_load_0_req_1); -- 
    cr_3920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => type_cast_1282_inst_req_1); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Sample/ra
      -- 
    ra_3794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_0, ack => zeropad3D_CP_2152_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Update/ca
      -- 
    ca_3799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_1, ack => zeropad3D_CP_2152_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/word_access_start/$exit
      -- CP-element group 119: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/word_access_start/word_0/$exit
      -- CP-element group 119: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/word_access_start/word_0/ra
      -- 
    ra_3816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1234_load_0_ack_0, ack => zeropad3D_CP_2152_elements(119)); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	116 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (12) 
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/word_access_complete/$exit
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/word_access_complete/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/word_access_complete/word_0/ca
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/LOAD_col_high_1234_Merge/$entry
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/LOAD_col_high_1234_Merge/$exit
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/LOAD_col_high_1234_Merge/merge_req
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/LOAD_col_high_1234_Merge/merge_ack
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Sample/rr
      -- 
    ca_3827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1234_load_0_ack_1, ack => zeropad3D_CP_2152_elements(120)); -- 
    rr_3840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(120), ack => type_cast_1238_inst_req_0); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Sample/ra
      -- 
    ra_3841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => zeropad3D_CP_2152_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	116 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Update/ca
      -- 
    ca_3846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => zeropad3D_CP_2152_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Sample/rr
      -- 
    rr_3854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(123), ack => type_cast_1258_inst_req_0); -- 
    zeropad3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(118) & zeropad3D_CP_2152_elements(122);
      gj_zeropad3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Sample/ra
      -- 
    ra_3855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1258_inst_ack_0, ack => zeropad3D_CP_2152_elements(124)); -- 
    -- CP-element group 125:  transition  input  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	116 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (6) 
      -- CP-element group 125: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Sample/rr
      -- 
    ca_3860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1258_inst_ack_1, ack => zeropad3D_CP_2152_elements(125)); -- 
    rr_3868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(125), ack => type_cast_1275_inst_req_0); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Sample/ra
      -- 
    ra_3869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1275_inst_ack_0, ack => zeropad3D_CP_2152_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	116 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	132 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Update/ca
      -- 
    ca_3874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1275_inst_ack_1, ack => zeropad3D_CP_2152_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	116 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (5) 
      -- CP-element group 128: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/word_access_start/$exit
      -- CP-element group 128: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/word_access_start/word_0/$exit
      -- CP-element group 128: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/word_access_start/word_0/ra
      -- 
    ra_3891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1278_load_0_ack_0, ack => zeropad3D_CP_2152_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	116 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (12) 
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/word_access_complete/$exit
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/word_access_complete/word_0/$exit
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/word_access_complete/word_0/ca
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/LOAD_row_high_1278_Merge/$entry
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/LOAD_row_high_1278_Merge/$exit
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/LOAD_row_high_1278_Merge/merge_req
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/LOAD_row_high_1278_Merge/merge_ack
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Sample/rr
      -- 
    ca_3902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1278_load_0_ack_1, ack => zeropad3D_CP_2152_elements(129)); -- 
    rr_3915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(129), ack => type_cast_1282_inst_req_0); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Sample/ra
      -- 
    ra_3916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1282_inst_ack_0, ack => zeropad3D_CP_2152_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	116 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Update/ca
      -- 
    ca_3921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1282_inst_ack_1, ack => zeropad3D_CP_2152_elements(131)); -- 
    -- CP-element group 132:  branch  join  transition  place  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	127 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (10) 
      -- CP-element group 132: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299__exit__
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300__entry__
      -- CP-element group 132: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/$exit
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300_dead_link/$entry
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300_eval_test/$entry
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300_eval_test/$exit
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300_eval_test/branch_req
      -- CP-element group 132: 	 branch_block_stmt_714/R_cmp176_1301_place
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300_if_link/$entry
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300_else_link/$entry
      -- 
    branch_req_3929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(132), ack => if_stmt_1300_branch_req_0); -- 
    zeropad3D_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(127) & zeropad3D_CP_2152_elements(131);
      gj_zeropad3D_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  fork  transition  place  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	824 
    -- CP-element group 133: 	825 
    -- CP-element group 133: 	827 
    -- CP-element group 133: 	828 
    -- CP-element group 133:  members (20) 
      -- CP-element group 133: 	 branch_block_stmt_714/if_stmt_1300_if_link/$exit
      -- CP-element group 133: 	 branch_block_stmt_714/if_stmt_1300_if_link/if_choice_transition
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/type_cast_1332/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/type_cast_1332/SplitProtocol/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/type_cast_1332/SplitProtocol/Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/type_cast_1332/SplitProtocol/Sample/rr
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/type_cast_1332/SplitProtocol/Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/type_cast_1332/SplitProtocol/Update/cr
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/type_cast_1336/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/type_cast_1336/SplitProtocol/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/type_cast_1336/SplitProtocol/Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/type_cast_1336/SplitProtocol/Sample/rr
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/type_cast_1336/SplitProtocol/Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/type_cast_1336/SplitProtocol/Update/cr
      -- 
    if_choice_transition_3934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1300_branch_ack_1, ack => zeropad3D_CP_2152_elements(133)); -- 
    rr_11332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => type_cast_1332_inst_req_0); -- 
    cr_11337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => type_cast_1332_inst_req_1); -- 
    rr_11355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => type_cast_1336_inst_req_0); -- 
    cr_11360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => type_cast_1336_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  place  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	801 
    -- CP-element group 134: 	802 
    -- CP-element group 134: 	804 
    -- CP-element group 134: 	805 
    -- CP-element group 134: 	806 
    -- CP-element group 134:  members (22) 
      -- CP-element group 134: 	 branch_block_stmt_714/if_stmt_1300_else_link/$exit
      -- CP-element group 134: 	 branch_block_stmt_714/if_stmt_1300_else_link/else_choice_transition
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Update/cr
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Update/cr
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1319/$entry
      -- 
    else_choice_transition_3938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1300_branch_ack_0, ack => zeropad3D_CP_2152_elements(134)); -- 
    cr_11201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(134), ack => type_cast_1318_inst_req_1); -- 
    rr_11196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(134), ack => type_cast_1318_inst_req_0); -- 
    cr_11232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(134), ack => type_cast_1310_inst_req_1); -- 
    rr_11227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(134), ack => type_cast_1310_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	833 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1340_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1340_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1340_Sample/ra
      -- 
    ra_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1340_inst_ack_0, ack => zeropad3D_CP_2152_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	833 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	149 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1340_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1340_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1340_Update/ca
      -- 
    ca_3957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1340_inst_ack_1, ack => zeropad3D_CP_2152_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	833 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (5) 
      -- CP-element group 137: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Sample/word_access_start/$exit
      -- CP-element group 137: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Sample/word_access_start/word_0/$exit
      -- CP-element group 137: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Sample/word_access_start/word_0/ra
      -- 
    ra_3974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1349_load_0_ack_0, ack => zeropad3D_CP_2152_elements(137)); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	833 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	147 
    -- CP-element group 138:  members (12) 
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Update/word_access_complete/$exit
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Update/word_access_complete/word_0/$exit
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Update/word_access_complete/word_0/ca
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Update/LOAD_pad_1349_Merge/$entry
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Update/LOAD_pad_1349_Merge/$exit
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Update/LOAD_pad_1349_Merge/merge_req
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Update/LOAD_pad_1349_Merge/merge_ack
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1419_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1419_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1419_Sample/rr
      -- 
    ca_3985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1349_load_0_ack_1, ack => zeropad3D_CP_2152_elements(138)); -- 
    rr_4145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(138), ack => type_cast_1419_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	833 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (5) 
      -- CP-element group 139: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Sample/word_access_start/$exit
      -- CP-element group 139: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Sample/word_access_start/word_0/$exit
      -- CP-element group 139: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Sample/word_access_start/word_0/ra
      -- 
    ra_4007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_1352_load_0_ack_0, ack => zeropad3D_CP_2152_elements(139)); -- 
    -- CP-element group 140:  transition  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	833 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	145 
    -- CP-element group 140:  members (12) 
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Update/word_access_complete/$exit
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Update/word_access_complete/word_0/$exit
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Update/word_access_complete/word_0/ca
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Update/LOAD_depth_high_1352_Merge/$entry
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Update/LOAD_depth_high_1352_Merge/$exit
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Update/LOAD_depth_high_1352_Merge/merge_req
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Update/LOAD_depth_high_1352_Merge/merge_ack
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1380_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1380_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1380_Sample/rr
      -- 
    ca_4018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_1352_load_0_ack_1, ack => zeropad3D_CP_2152_elements(140)); -- 
    rr_4131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(140), ack => type_cast_1380_inst_req_0); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	833 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (5) 
      -- CP-element group 141: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Sample/word_access_start/$exit
      -- CP-element group 141: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Sample/word_access_start/word_0/$exit
      -- CP-element group 141: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Sample/word_access_start/word_0/ra
      -- 
    ra_4057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1364_load_0_ack_0, ack => zeropad3D_CP_2152_elements(141)); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	833 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	149 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Update/word_access_complete/$exit
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Update/word_access_complete/word_0/$exit
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Update/word_access_complete/word_0/ca
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Update/ptr_deref_1364_Merge/$entry
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Update/ptr_deref_1364_Merge/$exit
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Update/ptr_deref_1364_Merge/merge_req
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Update/ptr_deref_1364_Merge/merge_ack
      -- 
    ca_4068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1364_load_0_ack_1, ack => zeropad3D_CP_2152_elements(142)); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	833 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (5) 
      -- CP-element group 143: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Sample/word_access_start/$exit
      -- CP-element group 143: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Sample/word_access_start/word_0/$exit
      -- CP-element group 143: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Sample/word_access_start/word_0/ra
      -- 
    ra_4107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1376_load_0_ack_0, ack => zeropad3D_CP_2152_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	833 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	149 
    -- CP-element group 144:  members (9) 
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Update/word_access_complete/$exit
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Update/word_access_complete/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Update/word_access_complete/word_0/ca
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Update/ptr_deref_1376_Merge/$entry
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Update/ptr_deref_1376_Merge/$exit
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Update/ptr_deref_1376_Merge/merge_req
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Update/ptr_deref_1376_Merge/merge_ack
      -- 
    ca_4118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1376_load_0_ack_1, ack => zeropad3D_CP_2152_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	140 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1380_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1380_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1380_Sample/ra
      -- 
    ra_4132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1380_inst_ack_0, ack => zeropad3D_CP_2152_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	833 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1380_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1380_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1380_Update/ca
      -- 
    ca_4137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1380_inst_ack_1, ack => zeropad3D_CP_2152_elements(146)); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	138 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1419_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1419_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1419_Sample/ra
      -- 
    ra_4146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1419_inst_ack_0, ack => zeropad3D_CP_2152_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	833 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1419_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1419_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1419_Update/ca
      -- 
    ca_4151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1419_inst_ack_1, ack => zeropad3D_CP_2152_elements(148)); -- 
    -- CP-element group 149:  join  fork  transition  place  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	136 
    -- CP-element group 149: 	142 
    -- CP-element group 149: 	144 
    -- CP-element group 149: 	146 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	844 
    -- CP-element group 149: 	845 
    -- CP-element group 149: 	847 
    -- CP-element group 149: 	848 
    -- CP-element group 149:  members (16) 
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244
      -- CP-element group 149: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461__exit__
      -- CP-element group 149: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/$exit
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/$entry
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/$entry
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/$entry
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/$entry
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/$entry
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Sample/rr
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Update/cr
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1470/$entry
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/$entry
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1477/$entry
      -- CP-element group 149: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/$entry
      -- 
    rr_11459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(149), ack => type_cast_1467_inst_req_0); -- 
    cr_11464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(149), ack => type_cast_1467_inst_req_1); -- 
    zeropad3D_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(136) & zeropad3D_CP_2152_elements(142) & zeropad3D_CP_2152_elements(144) & zeropad3D_CP_2152_elements(146) & zeropad3D_CP_2152_elements(148);
      gj_zeropad3D_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	854 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/type_cast_1488_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/type_cast_1488_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/type_cast_1488_Sample/ra
      -- 
    ra_4163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1488_inst_ack_0, ack => zeropad3D_CP_2152_elements(150)); -- 
    -- CP-element group 151:  branch  transition  place  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	854 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (13) 
      -- CP-element group 151: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496__exit__
      -- CP-element group 151: 	 branch_block_stmt_714/if_stmt_1497__entry__
      -- CP-element group 151: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/$exit
      -- CP-element group 151: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/type_cast_1488_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/type_cast_1488_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/type_cast_1488_Update/ca
      -- CP-element group 151: 	 branch_block_stmt_714/if_stmt_1497_dead_link/$entry
      -- CP-element group 151: 	 branch_block_stmt_714/if_stmt_1497_eval_test/$entry
      -- CP-element group 151: 	 branch_block_stmt_714/if_stmt_1497_eval_test/$exit
      -- CP-element group 151: 	 branch_block_stmt_714/if_stmt_1497_eval_test/branch_req
      -- CP-element group 151: 	 branch_block_stmt_714/R_cmp249_1498_place
      -- CP-element group 151: 	 branch_block_stmt_714/if_stmt_1497_if_link/$entry
      -- CP-element group 151: 	 branch_block_stmt_714/if_stmt_1497_else_link/$entry
      -- 
    ca_4168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1488_inst_ack_1, ack => zeropad3D_CP_2152_elements(151)); -- 
    branch_req_4176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(151), ack => if_stmt_1497_branch_req_0); -- 
    -- CP-element group 152:  transition  place  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	855 
    -- CP-element group 152:  members (5) 
      -- CP-element group 152: 	 branch_block_stmt_714/if_stmt_1497_if_link/$exit
      -- CP-element group 152: 	 branch_block_stmt_714/if_stmt_1497_if_link/if_choice_transition
      -- CP-element group 152: 	 branch_block_stmt_714/whilex_xbody244_ifx_xthen279
      -- CP-element group 152: 	 branch_block_stmt_714/whilex_xbody244_ifx_xthen279_PhiReq/$entry
      -- CP-element group 152: 	 branch_block_stmt_714/whilex_xbody244_ifx_xthen279_PhiReq/$exit
      -- 
    if_choice_transition_4181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1497_branch_ack_1, ack => zeropad3D_CP_2152_elements(152)); -- 
    -- CP-element group 153:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153: 	155 
    -- CP-element group 153: 	157 
    -- CP-element group 153:  members (27) 
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528__entry__
      -- CP-element group 153: 	 branch_block_stmt_714/merge_stmt_1503__exit__
      -- CP-element group 153: 	 branch_block_stmt_714/if_stmt_1497_else_link/$exit
      -- CP-element group 153: 	 branch_block_stmt_714/if_stmt_1497_else_link/else_choice_transition
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xbody244_lorx_xlhsx_xfalse251
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_update_start_
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_word_address_calculated
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_root_address_calculated
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Sample/word_access_start/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Sample/word_access_start/word_0/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Sample/word_access_start/word_0/rr
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Update/word_access_complete/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Update/word_access_complete/word_0/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Update/word_access_complete/word_0/cr
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/type_cast_1509_update_start_
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/type_cast_1509_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/type_cast_1509_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xbody244_lorx_xlhsx_xfalse251_PhiReq/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xbody244_lorx_xlhsx_xfalse251_PhiReq/$exit
      -- CP-element group 153: 	 branch_block_stmt_714/merge_stmt_1503_PhiReqMerge
      -- CP-element group 153: 	 branch_block_stmt_714/merge_stmt_1503_PhiAck/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/merge_stmt_1503_PhiAck/$exit
      -- CP-element group 153: 	 branch_block_stmt_714/merge_stmt_1503_PhiAck/dummy
      -- 
    else_choice_transition_4185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1497_branch_ack_0, ack => zeropad3D_CP_2152_elements(153)); -- 
    rr_4206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(153), ack => LOAD_row_high_1505_load_0_req_0); -- 
    cr_4217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(153), ack => LOAD_row_high_1505_load_0_req_1); -- 
    cr_4236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(153), ack => type_cast_1509_inst_req_1); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (5) 
      -- CP-element group 154: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Sample/word_access_start/$exit
      -- CP-element group 154: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Sample/word_access_start/word_0/$exit
      -- CP-element group 154: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Sample/word_access_start/word_0/ra
      -- 
    ra_4207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1505_load_0_ack_0, ack => zeropad3D_CP_2152_elements(154)); -- 
    -- CP-element group 155:  transition  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (12) 
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Update/word_access_complete/$exit
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Update/word_access_complete/word_0/$exit
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Update/word_access_complete/word_0/ca
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Update/LOAD_row_high_1505_Merge/$entry
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Update/LOAD_row_high_1505_Merge/$exit
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Update/LOAD_row_high_1505_Merge/merge_req
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/LOAD_row_high_1505_Update/LOAD_row_high_1505_Merge/merge_ack
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/type_cast_1509_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/type_cast_1509_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/type_cast_1509_Sample/rr
      -- 
    ca_4218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1505_load_0_ack_1, ack => zeropad3D_CP_2152_elements(155)); -- 
    rr_4231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(155), ack => type_cast_1509_inst_req_0); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/type_cast_1509_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/type_cast_1509_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/type_cast_1509_Sample/ra
      -- 
    ra_4232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1509_inst_ack_0, ack => zeropad3D_CP_2152_elements(156)); -- 
    -- CP-element group 157:  branch  transition  place  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	153 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (13) 
      -- CP-element group 157: 	 branch_block_stmt_714/if_stmt_1529__entry__
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528__exit__
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/$exit
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/type_cast_1509_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/type_cast_1509_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1506_to_assign_stmt_1528/type_cast_1509_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_714/if_stmt_1529_dead_link/$entry
      -- CP-element group 157: 	 branch_block_stmt_714/if_stmt_1529_eval_test/$entry
      -- CP-element group 157: 	 branch_block_stmt_714/if_stmt_1529_eval_test/$exit
      -- CP-element group 157: 	 branch_block_stmt_714/if_stmt_1529_eval_test/branch_req
      -- CP-element group 157: 	 branch_block_stmt_714/R_cmp260_1530_place
      -- CP-element group 157: 	 branch_block_stmt_714/if_stmt_1529_if_link/$entry
      -- CP-element group 157: 	 branch_block_stmt_714/if_stmt_1529_else_link/$entry
      -- 
    ca_4237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1509_inst_ack_1, ack => zeropad3D_CP_2152_elements(157)); -- 
    branch_req_4245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(157), ack => if_stmt_1529_branch_req_0); -- 
    -- CP-element group 158:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: 	161 
    -- CP-element group 158:  members (18) 
      -- CP-element group 158: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547__entry__
      -- CP-element group 158: 	 branch_block_stmt_714/merge_stmt_1535__exit__
      -- CP-element group 158: 	 branch_block_stmt_714/if_stmt_1529_if_link/$exit
      -- CP-element group 158: 	 branch_block_stmt_714/if_stmt_1529_if_link/if_choice_transition
      -- CP-element group 158: 	 branch_block_stmt_714/lorx_xlhsx_xfalse251_lorx_xlhsx_xfalse262
      -- CP-element group 158: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/$entry
      -- CP-element group 158: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/type_cast_1539_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/type_cast_1539_update_start_
      -- CP-element group 158: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/type_cast_1539_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/type_cast_1539_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/type_cast_1539_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/type_cast_1539_Update/cr
      -- CP-element group 158: 	 branch_block_stmt_714/lorx_xlhsx_xfalse251_lorx_xlhsx_xfalse262_PhiReq/$entry
      -- CP-element group 158: 	 branch_block_stmt_714/lorx_xlhsx_xfalse251_lorx_xlhsx_xfalse262_PhiReq/$exit
      -- CP-element group 158: 	 branch_block_stmt_714/merge_stmt_1535_PhiReqMerge
      -- CP-element group 158: 	 branch_block_stmt_714/merge_stmt_1535_PhiAck/$entry
      -- CP-element group 158: 	 branch_block_stmt_714/merge_stmt_1535_PhiAck/$exit
      -- CP-element group 158: 	 branch_block_stmt_714/merge_stmt_1535_PhiAck/dummy
      -- 
    if_choice_transition_4250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1529_branch_ack_1, ack => zeropad3D_CP_2152_elements(158)); -- 
    rr_4267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(158), ack => type_cast_1539_inst_req_0); -- 
    cr_4272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(158), ack => type_cast_1539_inst_req_1); -- 
    -- CP-element group 159:  transition  place  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	855 
    -- CP-element group 159:  members (5) 
      -- CP-element group 159: 	 branch_block_stmt_714/if_stmt_1529_else_link/$exit
      -- CP-element group 159: 	 branch_block_stmt_714/if_stmt_1529_else_link/else_choice_transition
      -- CP-element group 159: 	 branch_block_stmt_714/lorx_xlhsx_xfalse251_ifx_xthen279
      -- CP-element group 159: 	 branch_block_stmt_714/lorx_xlhsx_xfalse251_ifx_xthen279_PhiReq/$entry
      -- CP-element group 159: 	 branch_block_stmt_714/lorx_xlhsx_xfalse251_ifx_xthen279_PhiReq/$exit
      -- 
    else_choice_transition_4254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1529_branch_ack_0, ack => zeropad3D_CP_2152_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/type_cast_1539_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/type_cast_1539_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/type_cast_1539_Sample/ra
      -- 
    ra_4268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1539_inst_ack_0, ack => zeropad3D_CP_2152_elements(160)); -- 
    -- CP-element group 161:  branch  transition  place  input  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	158 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (13) 
      -- CP-element group 161: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547__exit__
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1548__entry__
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1548_else_link/$entry
      -- CP-element group 161: 	 branch_block_stmt_714/R_cmp267_1549_place
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1548_if_link/$entry
      -- CP-element group 161: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/$exit
      -- CP-element group 161: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/type_cast_1539_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/type_cast_1539_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_714/assign_stmt_1540_to_assign_stmt_1547/type_cast_1539_Update/ca
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1548_dead_link/$entry
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1548_eval_test/$entry
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1548_eval_test/$exit
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1548_eval_test/branch_req
      -- 
    ca_4273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1539_inst_ack_1, ack => zeropad3D_CP_2152_elements(161)); -- 
    branch_req_4281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(161), ack => if_stmt_1548_branch_req_0); -- 
    -- CP-element group 162:  transition  place  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	855 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_714/if_stmt_1548_if_link/if_choice_transition
      -- CP-element group 162: 	 branch_block_stmt_714/if_stmt_1548_if_link/$exit
      -- CP-element group 162: 	 branch_block_stmt_714/lorx_xlhsx_xfalse262_ifx_xthen279
      -- CP-element group 162: 	 branch_block_stmt_714/lorx_xlhsx_xfalse262_ifx_xthen279_PhiReq/$entry
      -- CP-element group 162: 	 branch_block_stmt_714/lorx_xlhsx_xfalse262_ifx_xthen279_PhiReq/$exit
      -- 
    if_choice_transition_4286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1548_branch_ack_1, ack => zeropad3D_CP_2152_elements(162)); -- 
    -- CP-element group 163:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163: 	165 
    -- CP-element group 163: 	167 
    -- CP-element group 163:  members (27) 
      -- CP-element group 163: 	 branch_block_stmt_714/merge_stmt_1554__exit__
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573__entry__
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/$entry
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/type_cast_1560_update_start_
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Update/word_access_complete/word_0/cr
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Update/word_access_complete/word_0/$entry
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Update/word_access_complete/$entry
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Sample/word_access_start/word_0/rr
      -- CP-element group 163: 	 branch_block_stmt_714/if_stmt_1548_else_link/else_choice_transition
      -- CP-element group 163: 	 branch_block_stmt_714/if_stmt_1548_else_link/$exit
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Sample/word_access_start/word_0/$entry
      -- CP-element group 163: 	 branch_block_stmt_714/lorx_xlhsx_xfalse262_lorx_xlhsx_xfalse269
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Sample/word_access_start/$entry
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_root_address_calculated
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_word_address_calculated
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_update_start_
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/type_cast_1560_Update/cr
      -- CP-element group 163: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/type_cast_1560_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_714/lorx_xlhsx_xfalse262_lorx_xlhsx_xfalse269_PhiReq/$entry
      -- CP-element group 163: 	 branch_block_stmt_714/lorx_xlhsx_xfalse262_lorx_xlhsx_xfalse269_PhiReq/$exit
      -- CP-element group 163: 	 branch_block_stmt_714/merge_stmt_1554_PhiReqMerge
      -- CP-element group 163: 	 branch_block_stmt_714/merge_stmt_1554_PhiAck/$entry
      -- CP-element group 163: 	 branch_block_stmt_714/merge_stmt_1554_PhiAck/$exit
      -- CP-element group 163: 	 branch_block_stmt_714/merge_stmt_1554_PhiAck/dummy
      -- 
    else_choice_transition_4290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1548_branch_ack_0, ack => zeropad3D_CP_2152_elements(163)); -- 
    cr_4322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(163), ack => LOAD_col_high_1556_load_0_req_1); -- 
    rr_4311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(163), ack => LOAD_col_high_1556_load_0_req_0); -- 
    cr_4341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(163), ack => type_cast_1560_inst_req_1); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Sample/word_access_start/word_0/ra
      -- CP-element group 164: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Sample/word_access_start/word_0/$exit
      -- CP-element group 164: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Sample/word_access_start/$exit
      -- CP-element group 164: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_sample_completed_
      -- 
    ra_4312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1556_load_0_ack_0, ack => zeropad3D_CP_2152_elements(164)); -- 
    -- CP-element group 165:  transition  input  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (12) 
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/type_cast_1560_Sample/rr
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/type_cast_1560_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Update/LOAD_col_high_1556_Merge/merge_ack
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Update/LOAD_col_high_1556_Merge/merge_req
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Update/LOAD_col_high_1556_Merge/$exit
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Update/LOAD_col_high_1556_Merge/$entry
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Update/word_access_complete/word_0/ca
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Update/word_access_complete/word_0/$exit
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Update/word_access_complete/$exit
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/LOAD_col_high_1556_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/type_cast_1560_Sample/$entry
      -- 
    ca_4323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1556_load_0_ack_1, ack => zeropad3D_CP_2152_elements(165)); -- 
    rr_4336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(165), ack => type_cast_1560_inst_req_0); -- 
    -- CP-element group 166:  transition  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/type_cast_1560_Sample/ra
      -- CP-element group 166: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/type_cast_1560_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/type_cast_1560_Sample/$exit
      -- 
    ra_4337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1560_inst_ack_0, ack => zeropad3D_CP_2152_elements(166)); -- 
    -- CP-element group 167:  branch  transition  place  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	163 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (13) 
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573__exit__
      -- CP-element group 167: 	 branch_block_stmt_714/if_stmt_1574__entry__
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/$exit
      -- CP-element group 167: 	 branch_block_stmt_714/R_cmp277_1575_place
      -- CP-element group 167: 	 branch_block_stmt_714/if_stmt_1574_else_link/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/if_stmt_1574_if_link/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/if_stmt_1574_eval_test/branch_req
      -- CP-element group 167: 	 branch_block_stmt_714/if_stmt_1574_eval_test/$exit
      -- CP-element group 167: 	 branch_block_stmt_714/if_stmt_1574_eval_test/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/if_stmt_1574_dead_link/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/type_cast_1560_Update/ca
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/type_cast_1560_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1557_to_assign_stmt_1573/type_cast_1560_update_completed_
      -- 
    ca_4342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1560_inst_ack_1, ack => zeropad3D_CP_2152_elements(167)); -- 
    branch_req_4350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(167), ack => if_stmt_1574_branch_req_0); -- 
    -- CP-element group 168:  fork  transition  place  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	167 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	184 
    -- CP-element group 168: 	185 
    -- CP-element group 168: 	187 
    -- CP-element group 168: 	189 
    -- CP-element group 168: 	191 
    -- CP-element group 168: 	193 
    -- CP-element group 168: 	195 
    -- CP-element group 168: 	197 
    -- CP-element group 168: 	199 
    -- CP-element group 168: 	202 
    -- CP-element group 168:  members (46) 
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743__entry__
      -- CP-element group 168: 	 branch_block_stmt_714/merge_stmt_1638__exit__
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1738_update_start_
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_update_start_
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1713_complete/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1731_Update/cr
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1706_update_start_
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Update/word_access_complete/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1731_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/lorx_xlhsx_xfalse269_ifx_xelse300
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1642_Update/cr
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1642_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1731_update_start_
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1642_Sample/rr
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_update_start_
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1642_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_final_index_sum_regn_Update/req
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1642_update_start_
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1642_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1738_complete/req
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_final_index_sum_regn_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Update/word_access_complete/word_0/cr
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Update/word_access_complete/word_0/cr
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Update/word_access_complete/word_0/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1738_complete/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Update/word_access_complete/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_final_index_sum_regn_update_start
      -- CP-element group 168: 	 branch_block_stmt_714/if_stmt_1574_if_link/if_choice_transition
      -- CP-element group 168: 	 branch_block_stmt_714/if_stmt_1574_if_link/$exit
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_final_index_sum_regn_Update/req
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1713_update_start_
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_final_index_sum_regn_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1706_Update/cr
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_final_index_sum_regn_update_start
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Update/word_access_complete/word_0/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1713_complete/req
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1706_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/lorx_xlhsx_xfalse269_ifx_xelse300_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/lorx_xlhsx_xfalse269_ifx_xelse300_PhiReq/$exit
      -- CP-element group 168: 	 branch_block_stmt_714/merge_stmt_1638_PhiReqMerge
      -- CP-element group 168: 	 branch_block_stmt_714/merge_stmt_1638_PhiAck/$entry
      -- CP-element group 168: 	 branch_block_stmt_714/merge_stmt_1638_PhiAck/$exit
      -- CP-element group 168: 	 branch_block_stmt_714/merge_stmt_1638_PhiAck/dummy
      -- 
    if_choice_transition_4355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1574_branch_ack_1, ack => zeropad3D_CP_2152_elements(168)); -- 
    cr_4642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(168), ack => type_cast_1731_inst_req_1); -- 
    cr_4518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(168), ack => type_cast_1642_inst_req_1); -- 
    rr_4513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(168), ack => type_cast_1642_inst_req_0); -- 
    req_4563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(168), ack => array_obj_ref_1712_index_offset_req_1); -- 
    req_4688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(168), ack => addr_of_1738_final_reg_req_1); -- 
    cr_4738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(168), ack => ptr_deref_1741_store_0_req_1); -- 
    cr_4623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(168), ack => ptr_deref_1717_load_0_req_1); -- 
    req_4673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(168), ack => array_obj_ref_1737_index_offset_req_1); -- 
    cr_4532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(168), ack => type_cast_1706_inst_req_1); -- 
    req_4578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(168), ack => addr_of_1713_final_reg_req_1); -- 
    -- CP-element group 169:  transition  place  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	855 
    -- CP-element group 169:  members (5) 
      -- CP-element group 169: 	 branch_block_stmt_714/lorx_xlhsx_xfalse269_ifx_xthen279
      -- CP-element group 169: 	 branch_block_stmt_714/if_stmt_1574_else_link/else_choice_transition
      -- CP-element group 169: 	 branch_block_stmt_714/if_stmt_1574_else_link/$exit
      -- CP-element group 169: 	 branch_block_stmt_714/lorx_xlhsx_xfalse269_ifx_xthen279_PhiReq/$entry
      -- CP-element group 169: 	 branch_block_stmt_714/lorx_xlhsx_xfalse269_ifx_xthen279_PhiReq/$exit
      -- 
    else_choice_transition_4359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1574_branch_ack_0, ack => zeropad3D_CP_2152_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	855 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1584_Sample/ra
      -- CP-element group 170: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1584_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1584_sample_completed_
      -- 
    ra_4373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1584_inst_ack_0, ack => zeropad3D_CP_2152_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	855 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	174 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1584_Update/ca
      -- CP-element group 171: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1584_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1584_update_completed_
      -- 
    ca_4378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1584_inst_ack_1, ack => zeropad3D_CP_2152_elements(171)); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	855 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1589_Sample/ra
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1589_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1589_sample_completed_
      -- 
    ra_4387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1589_inst_ack_0, ack => zeropad3D_CP_2152_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	855 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1589_Update/ca
      -- CP-element group 173: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1589_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1589_update_completed_
      -- 
    ca_4392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1589_inst_ack_1, ack => zeropad3D_CP_2152_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	171 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1623_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1623_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1623_sample_start_
      -- 
    rr_4400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(174), ack => type_cast_1623_inst_req_0); -- 
    zeropad3D_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(171) & zeropad3D_CP_2152_elements(173);
      gj_zeropad3D_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1623_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1623_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1623_sample_completed_
      -- 
    ra_4401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1623_inst_ack_0, ack => zeropad3D_CP_2152_elements(175)); -- 
    -- CP-element group 176:  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	855 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (16) 
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_final_index_sum_regn_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_index_scale_1/scale_rename_ack
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_index_scale_1/scale_rename_req
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_index_scale_1/$exit
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_index_scale_1/$entry
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_index_resize_1/index_resize_ack
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_index_resize_1/index_resize_req
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_index_resize_1/$exit
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_index_resize_1/$entry
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_index_computed_1
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_index_scaled_1
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_index_resized_1
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1623_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1623_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1623_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_final_index_sum_regn_Sample/req
      -- 
    ca_4406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1623_inst_ack_1, ack => zeropad3D_CP_2152_elements(176)); -- 
    req_4431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(176), ack => array_obj_ref_1629_index_offset_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	183 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_final_index_sum_regn_sample_complete
      -- CP-element group 177: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_final_index_sum_regn_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_final_index_sum_regn_Sample/ack
      -- 
    ack_4432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1629_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(177)); -- 
    -- CP-element group 178:  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	855 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (11) 
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_offset_calculated
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_root_address_calculated
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/addr_of_1630_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/addr_of_1630_request/req
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/addr_of_1630_request/$entry
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_base_plus_offset/sum_rename_ack
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_base_plus_offset/sum_rename_req
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_base_plus_offset/$exit
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_base_plus_offset/$entry
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_final_index_sum_regn_Update/ack
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_final_index_sum_regn_Update/$exit
      -- 
    ack_4437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1629_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(178)); -- 
    req_4446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(178), ack => addr_of_1630_final_reg_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/addr_of_1630_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/addr_of_1630_request/ack
      -- CP-element group 179: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/addr_of_1630_request/$exit
      -- 
    ack_4447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1630_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(179)); -- 
    -- CP-element group 180:  join  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	855 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (28) 
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_base_plus_offset/sum_rename_req
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_base_plus_offset/$exit
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_base_plus_offset/sum_rename_ack
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_base_plus_offset/$entry
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_base_addr_resize/base_resize_ack
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_base_addr_resize/base_resize_req
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_base_addr_resize/$exit
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_base_addr_resize/$entry
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_base_address_resized
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_root_address_calculated
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_word_address_calculated
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_base_address_calculated
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/addr_of_1630_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/addr_of_1630_complete/ack
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/addr_of_1630_complete/$exit
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Sample/word_access_start/word_0/rr
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Sample/word_access_start/word_0/$entry
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Sample/word_access_start/$entry
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Sample/ptr_deref_1633_Split/split_ack
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Sample/ptr_deref_1633_Split/split_req
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Sample/ptr_deref_1633_Split/$exit
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Sample/ptr_deref_1633_Split/$entry
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_word_addrgen/root_register_ack
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_word_addrgen/root_register_req
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_word_addrgen/$exit
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_word_addrgen/$entry
      -- 
    ack_4452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1630_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(180)); -- 
    rr_4490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(180), ack => ptr_deref_1633_store_0_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (5) 
      -- CP-element group 181: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Sample/word_access_start/word_0/ra
      -- CP-element group 181: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Sample/word_access_start/word_0/$exit
      -- CP-element group 181: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Sample/word_access_start/$exit
      -- CP-element group 181: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Sample/$exit
      -- 
    ra_4491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1633_store_0_ack_0, ack => zeropad3D_CP_2152_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	855 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (5) 
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Update/word_access_complete/word_0/ca
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Update/word_access_complete/word_0/$exit
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Update/word_access_complete/$exit
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Update/$exit
      -- 
    ca_4502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1633_store_0_ack_1, ack => zeropad3D_CP_2152_elements(182)); -- 
    -- CP-element group 183:  join  transition  place  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	177 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	856 
    -- CP-element group 183:  members (5) 
      -- CP-element group 183: 	 branch_block_stmt_714/ifx_xthen279_ifx_xend348
      -- CP-element group 183: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636__exit__
      -- CP-element group 183: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/$exit
      -- CP-element group 183: 	 branch_block_stmt_714/ifx_xthen279_ifx_xend348_PhiReq/$entry
      -- CP-element group 183: 	 branch_block_stmt_714/ifx_xthen279_ifx_xend348_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(177) & zeropad3D_CP_2152_elements(182);
      gj_zeropad3D_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	168 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1642_Sample/ra
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1642_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1642_sample_completed_
      -- 
    ra_4514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1642_inst_ack_0, ack => zeropad3D_CP_2152_elements(184)); -- 
    -- CP-element group 185:  fork  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	168 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185: 	194 
    -- CP-element group 185:  members (9) 
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1706_Sample/rr
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1706_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1731_Sample/rr
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1706_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1731_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1642_Update/ca
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1642_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1731_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1642_update_completed_
      -- 
    ca_4519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1642_inst_ack_1, ack => zeropad3D_CP_2152_elements(185)); -- 
    rr_4527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(185), ack => type_cast_1706_inst_req_0); -- 
    rr_4637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(185), ack => type_cast_1731_inst_req_0); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1706_Sample/ra
      -- CP-element group 186: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1706_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1706_sample_completed_
      -- 
    ra_4528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1706_inst_ack_0, ack => zeropad3D_CP_2152_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	168 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (16) 
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1706_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_final_index_sum_regn_Sample/req
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_final_index_sum_regn_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_index_scale_1/scale_rename_ack
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_index_scale_1/scale_rename_req
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_index_scale_1/$exit
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_index_scale_1/$entry
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_index_resize_1/index_resize_ack
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_index_resize_1/index_resize_req
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_index_resize_1/$exit
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_index_resize_1/$entry
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_index_computed_1
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_index_scaled_1
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_index_resized_1
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1706_Update/ca
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1706_Update/$exit
      -- 
    ca_4533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1706_inst_ack_1, ack => zeropad3D_CP_2152_elements(187)); -- 
    req_4558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(187), ack => array_obj_ref_1712_index_offset_req_0); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	203 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_final_index_sum_regn_Sample/ack
      -- CP-element group 188: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_final_index_sum_regn_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_final_index_sum_regn_sample_complete
      -- 
    ack_4559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1712_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	168 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (11) 
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1713_request/req
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1713_request/$entry
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_base_plus_offset/sum_rename_ack
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_base_plus_offset/sum_rename_req
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_base_plus_offset/$exit
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_base_plus_offset/$entry
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_final_index_sum_regn_Update/ack
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_final_index_sum_regn_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_offset_calculated
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1712_root_address_calculated
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1713_sample_start_
      -- 
    ack_4564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1712_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(189)); -- 
    req_4573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(189), ack => addr_of_1713_final_reg_req_0); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1713_request/ack
      -- CP-element group 190: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1713_request/$exit
      -- CP-element group 190: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1713_sample_completed_
      -- 
    ack_4574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1713_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(190)); -- 
    -- CP-element group 191:  join  fork  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	168 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (24) 
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_base_addr_resize/$entry
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1713_complete/$exit
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_base_addr_resize/$exit
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_base_address_resized
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_root_address_calculated
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_word_address_calculated
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_base_address_calculated
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Sample/word_access_start/word_0/rr
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Sample/word_access_start/word_0/$entry
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1713_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Sample/word_access_start/$entry
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_word_addrgen/root_register_ack
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_word_addrgen/root_register_req
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_word_addrgen/$exit
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_word_addrgen/$entry
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_base_plus_offset/sum_rename_ack
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_base_plus_offset/sum_rename_req
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_base_plus_offset/$exit
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1713_complete/ack
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_base_plus_offset/$entry
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_base_addr_resize/base_resize_ack
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_base_addr_resize/base_resize_req
      -- 
    ack_4579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1713_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(191)); -- 
    rr_4612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(191), ack => ptr_deref_1717_load_0_req_0); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (5) 
      -- CP-element group 192: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Sample/word_access_start/word_0/ra
      -- CP-element group 192: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Sample/word_access_start/word_0/$exit
      -- CP-element group 192: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Sample/word_access_start/$exit
      -- CP-element group 192: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Sample/$exit
      -- 
    ra_4613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_load_0_ack_0, ack => zeropad3D_CP_2152_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	168 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	200 
    -- CP-element group 193:  members (9) 
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Update/ptr_deref_1717_Merge/merge_ack
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Update/ptr_deref_1717_Merge/merge_req
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Update/ptr_deref_1717_Merge/$exit
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Update/ptr_deref_1717_Merge/$entry
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Update/word_access_complete/word_0/ca
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Update/word_access_complete/word_0/$exit
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Update/word_access_complete/$exit
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1717_update_completed_
      -- 
    ca_4624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_load_0_ack_1, ack => zeropad3D_CP_2152_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	185 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1731_Sample/ra
      -- CP-element group 194: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1731_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1731_sample_completed_
      -- 
    ra_4638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1731_inst_ack_0, ack => zeropad3D_CP_2152_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	168 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (16) 
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_index_scale_1/scale_rename_ack
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_index_scale_1/scale_rename_req
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1731_Update/ca
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1731_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_index_scale_1/$exit
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_index_scale_1/$entry
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/type_cast_1731_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_index_resize_1/index_resize_ack
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_index_resize_1/index_resize_req
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_index_resize_1/$exit
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_index_resize_1/$entry
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_index_computed_1
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_final_index_sum_regn_Sample/req
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_final_index_sum_regn_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_index_scaled_1
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_index_resized_1
      -- 
    ca_4643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1731_inst_ack_1, ack => zeropad3D_CP_2152_elements(195)); -- 
    req_4668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(195), ack => array_obj_ref_1737_index_offset_req_0); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	203 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_final_index_sum_regn_Sample/ack
      -- CP-element group 196: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_final_index_sum_regn_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_final_index_sum_regn_sample_complete
      -- 
    ack_4669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1737_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	168 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (11) 
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1738_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1738_request/req
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_base_plus_offset/sum_rename_ack
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_base_plus_offset/sum_rename_req
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_base_plus_offset/$exit
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_base_plus_offset/$entry
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_final_index_sum_regn_Update/ack
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_final_index_sum_regn_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1738_request/$entry
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_offset_calculated
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/array_obj_ref_1737_root_address_calculated
      -- 
    ack_4674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1737_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(197)); -- 
    req_4683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(197), ack => addr_of_1738_final_reg_req_0); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1738_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1738_request/ack
      -- CP-element group 198: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1738_request/$exit
      -- 
    ack_4684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1738_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(198)); -- 
    -- CP-element group 199:  fork  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	168 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (19) 
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_base_addr_resize/$exit
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1738_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_base_addr_resize/$entry
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_base_address_resized
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_word_addrgen/root_register_ack
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_root_address_calculated
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_word_address_calculated
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_word_addrgen/root_register_req
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_word_addrgen/$exit
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_base_address_calculated
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_word_addrgen/$entry
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1738_complete/ack
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_base_plus_offset/sum_rename_ack
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/addr_of_1738_complete/$exit
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_base_plus_offset/sum_rename_req
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_base_plus_offset/$exit
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_base_plus_offset/$entry
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_base_addr_resize/base_resize_ack
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_base_addr_resize/base_resize_req
      -- 
    ack_4689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1738_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	193 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (9) 
      -- CP-element group 200: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Sample/ptr_deref_1741_Split/$exit
      -- CP-element group 200: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Sample/word_access_start/word_0/rr
      -- CP-element group 200: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Sample/ptr_deref_1741_Split/$entry
      -- CP-element group 200: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Sample/word_access_start/word_0/$entry
      -- CP-element group 200: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Sample/word_access_start/$entry
      -- CP-element group 200: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Sample/ptr_deref_1741_Split/split_ack
      -- CP-element group 200: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Sample/ptr_deref_1741_Split/split_req
      -- 
    rr_4727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(200), ack => ptr_deref_1741_store_0_req_0); -- 
    zeropad3D_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(193) & zeropad3D_CP_2152_elements(199);
      gj_zeropad3D_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (5) 
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Sample/word_access_start/word_0/ra
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Sample/word_access_start/word_0/$exit
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Sample/word_access_start/$exit
      -- 
    ra_4728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1741_store_0_ack_0, ack => zeropad3D_CP_2152_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	168 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (5) 
      -- CP-element group 202: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Update/word_access_complete/$exit
      -- CP-element group 202: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Update/word_access_complete/word_0/ca
      -- CP-element group 202: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/ptr_deref_1741_Update/word_access_complete/word_0/$exit
      -- 
    ca_4739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1741_store_0_ack_1, ack => zeropad3D_CP_2152_elements(202)); -- 
    -- CP-element group 203:  join  transition  place  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	188 
    -- CP-element group 203: 	196 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	856 
    -- CP-element group 203:  members (5) 
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743__exit__
      -- CP-element group 203: 	 branch_block_stmt_714/ifx_xelse300_ifx_xend348
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1643_to_assign_stmt_1743/$exit
      -- CP-element group 203: 	 branch_block_stmt_714/ifx_xelse300_ifx_xend348_PhiReq/$entry
      -- CP-element group 203: 	 branch_block_stmt_714/ifx_xelse300_ifx_xend348_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(188) & zeropad3D_CP_2152_elements(196) & zeropad3D_CP_2152_elements(202);
      gj_zeropad3D_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	856 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/type_cast_1749_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/type_cast_1749_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/type_cast_1749_Sample/ra
      -- 
    ra_4751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1749_inst_ack_0, ack => zeropad3D_CP_2152_elements(204)); -- 
    -- CP-element group 205:  branch  transition  place  input  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	856 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205: 	207 
    -- CP-element group 205:  members (13) 
      -- CP-element group 205: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763__exit__
      -- CP-element group 205: 	 branch_block_stmt_714/if_stmt_1764__entry__
      -- CP-element group 205: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/$exit
      -- CP-element group 205: 	 branch_block_stmt_714/R_cmp356_1765_place
      -- CP-element group 205: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/type_cast_1749_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/type_cast_1749_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/type_cast_1749_Update/ca
      -- CP-element group 205: 	 branch_block_stmt_714/if_stmt_1764_dead_link/$entry
      -- CP-element group 205: 	 branch_block_stmt_714/if_stmt_1764_eval_test/$entry
      -- CP-element group 205: 	 branch_block_stmt_714/if_stmt_1764_eval_test/$exit
      -- CP-element group 205: 	 branch_block_stmt_714/if_stmt_1764_eval_test/branch_req
      -- CP-element group 205: 	 branch_block_stmt_714/if_stmt_1764_if_link/$entry
      -- CP-element group 205: 	 branch_block_stmt_714/if_stmt_1764_else_link/$entry
      -- 
    ca_4756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1749_inst_ack_1, ack => zeropad3D_CP_2152_elements(205)); -- 
    branch_req_4764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(205), ack => if_stmt_1764_branch_req_0); -- 
    -- CP-element group 206:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	865 
    -- CP-element group 206: 	866 
    -- CP-element group 206: 	868 
    -- CP-element group 206: 	869 
    -- CP-element group 206: 	871 
    -- CP-element group 206: 	872 
    -- CP-element group 206:  members (40) 
      -- CP-element group 206: 	 branch_block_stmt_714/merge_stmt_1770__exit__
      -- CP-element group 206: 	 branch_block_stmt_714/assign_stmt_1776__entry__
      -- CP-element group 206: 	 branch_block_stmt_714/assign_stmt_1776__exit__
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xend348_ifx_xthen358
      -- CP-element group 206: 	 branch_block_stmt_714/if_stmt_1764_if_link/$exit
      -- CP-element group 206: 	 branch_block_stmt_714/if_stmt_1764_if_link/if_choice_transition
      -- CP-element group 206: 	 branch_block_stmt_714/assign_stmt_1776/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/assign_stmt_1776/$exit
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xend348_ifx_xthen358_PhiReq/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xend348_ifx_xthen358_PhiReq/$exit
      -- CP-element group 206: 	 branch_block_stmt_714/merge_stmt_1770_PhiReqMerge
      -- CP-element group 206: 	 branch_block_stmt_714/merge_stmt_1770_PhiAck/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/merge_stmt_1770_PhiAck/$exit
      -- CP-element group 206: 	 branch_block_stmt_714/merge_stmt_1770_PhiAck/dummy
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/type_cast_1872/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/type_cast_1872/SplitProtocol/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/type_cast_1872/SplitProtocol/Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/type_cast_1872/SplitProtocol/Sample/rr
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/type_cast_1872/SplitProtocol/Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/type_cast_1872/SplitProtocol/Update/cr
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1866/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1866/SplitProtocol/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1866/SplitProtocol/Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1866/SplitProtocol/Sample/rr
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1866/SplitProtocol/Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1866/SplitProtocol/Update/cr
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1860/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1860/SplitProtocol/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1860/SplitProtocol/Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1860/SplitProtocol/Sample/rr
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1860/SplitProtocol/Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1860/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1764_branch_ack_1, ack => zeropad3D_CP_2152_elements(206)); -- 
    rr_11665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(206), ack => type_cast_1872_inst_req_0); -- 
    cr_11670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(206), ack => type_cast_1872_inst_req_1); -- 
    rr_11688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(206), ack => type_cast_1866_inst_req_0); -- 
    cr_11693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(206), ack => type_cast_1866_inst_req_1); -- 
    rr_11711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(206), ack => type_cast_1860_inst_req_0); -- 
    cr_11716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(206), ack => type_cast_1860_inst_req_1); -- 
    -- CP-element group 207:  fork  transition  place  input  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	205 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207: 	209 
    -- CP-element group 207: 	210 
    -- CP-element group 207: 	211 
    -- CP-element group 207: 	213 
    -- CP-element group 207: 	216 
    -- CP-element group 207: 	218 
    -- CP-element group 207: 	219 
    -- CP-element group 207: 	220 
    -- CP-element group 207: 	222 
    -- CP-element group 207:  members (54) 
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849__entry__
      -- CP-element group 207: 	 branch_block_stmt_714/merge_stmt_1778__exit__
      -- CP-element group 207: 	 branch_block_stmt_714/ifx_xend348_ifx_xelse363
      -- CP-element group 207: 	 branch_block_stmt_714/if_stmt_1764_else_link/$exit
      -- CP-element group 207: 	 branch_block_stmt_714/if_stmt_1764_else_link/else_choice_transition
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1788_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1788_update_start_
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1788_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1788_Sample/rr
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1788_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1788_Update/cr
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_update_start_
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_word_address_calculated
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_root_address_calculated
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Sample/word_access_start/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Sample/word_access_start/word_0/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Sample/word_access_start/word_0/rr
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Update/word_access_complete/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Update/word_access_complete/word_0/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Update/word_access_complete/word_0/cr
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1795_update_start_
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1795_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1795_Update/cr
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1809_update_start_
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1809_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1809_Update/cr
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1825_update_start_
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1825_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1825_Update/cr
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_update_start_
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_word_address_calculated
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_root_address_calculated
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Sample/word_access_start/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Sample/word_access_start/word_0/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Sample/word_access_start/word_0/rr
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Update/word_access_complete/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Update/word_access_complete/word_0/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Update/word_access_complete/word_0/cr
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1832_update_start_
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1832_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1832_Update/cr
      -- CP-element group 207: 	 branch_block_stmt_714/ifx_xend348_ifx_xelse363_PhiReq/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/ifx_xend348_ifx_xelse363_PhiReq/$exit
      -- CP-element group 207: 	 branch_block_stmt_714/merge_stmt_1778_PhiReqMerge
      -- CP-element group 207: 	 branch_block_stmt_714/merge_stmt_1778_PhiAck/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/merge_stmt_1778_PhiAck/$exit
      -- CP-element group 207: 	 branch_block_stmt_714/merge_stmt_1778_PhiAck/dummy
      -- 
    else_choice_transition_4773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1764_branch_ack_0, ack => zeropad3D_CP_2152_elements(207)); -- 
    rr_4789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(207), ack => type_cast_1788_inst_req_0); -- 
    cr_4794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(207), ack => type_cast_1788_inst_req_1); -- 
    rr_4811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(207), ack => LOAD_col_high_1791_load_0_req_0); -- 
    cr_4822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(207), ack => LOAD_col_high_1791_load_0_req_1); -- 
    cr_4841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(207), ack => type_cast_1795_inst_req_1); -- 
    cr_4855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(207), ack => type_cast_1809_inst_req_1); -- 
    cr_4869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(207), ack => type_cast_1825_inst_req_1); -- 
    rr_4886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(207), ack => LOAD_row_high_1828_load_0_req_0); -- 
    cr_4897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(207), ack => LOAD_row_high_1828_load_0_req_1); -- 
    cr_4916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(207), ack => type_cast_1832_inst_req_1); -- 
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1788_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1788_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1788_Sample/ra
      -- 
    ra_4790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1788_inst_ack_0, ack => zeropad3D_CP_2152_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	214 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1788_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1788_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1788_Update/ca
      -- 
    ca_4795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1788_inst_ack_1, ack => zeropad3D_CP_2152_elements(209)); -- 
    -- CP-element group 210:  transition  input  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	207 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (5) 
      -- CP-element group 210: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_sample_completed_
      -- CP-element group 210: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Sample/$exit
      -- CP-element group 210: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Sample/word_access_start/$exit
      -- CP-element group 210: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Sample/word_access_start/word_0/$exit
      -- CP-element group 210: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Sample/word_access_start/word_0/ra
      -- 
    ra_4812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1791_load_0_ack_0, ack => zeropad3D_CP_2152_elements(210)); -- 
    -- CP-element group 211:  transition  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	207 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	212 
    -- CP-element group 211:  members (12) 
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_update_completed_
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Update/$exit
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Update/word_access_complete/$exit
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Update/word_access_complete/word_0/$exit
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Update/word_access_complete/word_0/ca
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Update/LOAD_col_high_1791_Merge/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Update/LOAD_col_high_1791_Merge/$exit
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Update/LOAD_col_high_1791_Merge/merge_req
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_col_high_1791_Update/LOAD_col_high_1791_Merge/merge_ack
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1795_sample_start_
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1795_Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1795_Sample/rr
      -- 
    ca_4823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1791_load_0_ack_1, ack => zeropad3D_CP_2152_elements(211)); -- 
    rr_4836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(211), ack => type_cast_1795_inst_req_0); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	211 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1795_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1795_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1795_Sample/ra
      -- 
    ra_4837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1795_inst_ack_0, ack => zeropad3D_CP_2152_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	207 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1795_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1795_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1795_Update/ca
      -- 
    ca_4842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1795_inst_ack_1, ack => zeropad3D_CP_2152_elements(213)); -- 
    -- CP-element group 214:  join  transition  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	209 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1809_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1809_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1809_Sample/rr
      -- 
    rr_4850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(214), ack => type_cast_1809_inst_req_0); -- 
    zeropad3D_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(209) & zeropad3D_CP_2152_elements(213);
      gj_zeropad3D_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1809_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1809_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1809_Sample/ra
      -- 
    ra_4851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1809_inst_ack_0, ack => zeropad3D_CP_2152_elements(215)); -- 
    -- CP-element group 216:  transition  input  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	207 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (6) 
      -- CP-element group 216: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1809_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1809_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1809_Update/ca
      -- CP-element group 216: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1825_sample_start_
      -- CP-element group 216: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1825_Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1825_Sample/rr
      -- 
    ca_4856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1809_inst_ack_1, ack => zeropad3D_CP_2152_elements(216)); -- 
    rr_4864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(216), ack => type_cast_1825_inst_req_0); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1825_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1825_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1825_Sample/ra
      -- 
    ra_4865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1825_inst_ack_0, ack => zeropad3D_CP_2152_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	207 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	223 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1825_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1825_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1825_Update/ca
      -- 
    ca_4870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1825_inst_ack_1, ack => zeropad3D_CP_2152_elements(218)); -- 
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	207 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Sample/word_access_start/$exit
      -- CP-element group 219: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Sample/word_access_start/word_0/$exit
      -- CP-element group 219: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Sample/word_access_start/word_0/ra
      -- 
    ra_4887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1828_load_0_ack_0, ack => zeropad3D_CP_2152_elements(219)); -- 
    -- CP-element group 220:  transition  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	207 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220:  members (12) 
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Update/word_access_complete/$exit
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Update/word_access_complete/word_0/$exit
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Update/word_access_complete/word_0/ca
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Update/LOAD_row_high_1828_Merge/$entry
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Update/LOAD_row_high_1828_Merge/$exit
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Update/LOAD_row_high_1828_Merge/merge_req
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/LOAD_row_high_1828_Update/LOAD_row_high_1828_Merge/merge_ack
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1832_sample_start_
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1832_Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1832_Sample/rr
      -- 
    ca_4898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1828_load_0_ack_1, ack => zeropad3D_CP_2152_elements(220)); -- 
    rr_4911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(220), ack => type_cast_1832_inst_req_0); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1832_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1832_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1832_Sample/ra
      -- 
    ra_4912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1832_inst_ack_0, ack => zeropad3D_CP_2152_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	207 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1832_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1832_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/type_cast_1832_Update/ca
      -- 
    ca_4917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1832_inst_ack_1, ack => zeropad3D_CP_2152_elements(222)); -- 
    -- CP-element group 223:  branch  join  transition  place  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	218 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (10) 
      -- CP-element group 223: 	 branch_block_stmt_714/if_stmt_1850__entry__
      -- CP-element group 223: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849__exit__
      -- CP-element group 223: 	 branch_block_stmt_714/assign_stmt_1784_to_assign_stmt_1849/$exit
      -- CP-element group 223: 	 branch_block_stmt_714/if_stmt_1850_dead_link/$entry
      -- CP-element group 223: 	 branch_block_stmt_714/if_stmt_1850_eval_test/$entry
      -- CP-element group 223: 	 branch_block_stmt_714/if_stmt_1850_eval_test/$exit
      -- CP-element group 223: 	 branch_block_stmt_714/if_stmt_1850_eval_test/branch_req
      -- CP-element group 223: 	 branch_block_stmt_714/R_cmp390_1851_place
      -- CP-element group 223: 	 branch_block_stmt_714/if_stmt_1850_if_link/$entry
      -- CP-element group 223: 	 branch_block_stmt_714/if_stmt_1850_else_link/$entry
      -- 
    branch_req_4925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(223), ack => if_stmt_1850_branch_req_0); -- 
    zeropad3D_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(218) & zeropad3D_CP_2152_elements(222);
      gj_zeropad3D_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  place  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	880 
    -- CP-element group 224: 	881 
    -- CP-element group 224: 	883 
    -- CP-element group 224: 	884 
    -- CP-element group 224:  members (20) 
      -- CP-element group 224: 	 branch_block_stmt_714/if_stmt_1850_if_link/$exit
      -- CP-element group 224: 	 branch_block_stmt_714/if_stmt_1850_if_link/if_choice_transition
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/type_cast_1886/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/type_cast_1886/SplitProtocol/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/type_cast_1886/SplitProtocol/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/type_cast_1886/SplitProtocol/Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/type_cast_1886/SplitProtocol/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/type_cast_1886/SplitProtocol/Update/cr
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/type_cast_1882/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/type_cast_1882/SplitProtocol/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/type_cast_1882/SplitProtocol/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/type_cast_1882/SplitProtocol/Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/type_cast_1882/SplitProtocol/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/type_cast_1882/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1850_branch_ack_1, ack => zeropad3D_CP_2152_elements(224)); -- 
    rr_11744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(224), ack => type_cast_1886_inst_req_0); -- 
    cr_11749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(224), ack => type_cast_1886_inst_req_1); -- 
    rr_11767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(224), ack => type_cast_1882_inst_req_0); -- 
    cr_11772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(224), ack => type_cast_1882_inst_req_1); -- 
    -- CP-element group 225:  fork  transition  place  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	857 
    -- CP-element group 225: 	858 
    -- CP-element group 225: 	859 
    -- CP-element group 225: 	861 
    -- CP-element group 225: 	862 
    -- CP-element group 225:  members (22) 
      -- CP-element group 225: 	 branch_block_stmt_714/if_stmt_1850_else_link/$exit
      -- CP-element group 225: 	 branch_block_stmt_714/if_stmt_1850_else_link/else_choice_transition
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1869/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1868/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1868/SplitProtocol/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1868/SplitProtocol/Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1868/SplitProtocol/Sample/rr
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1868/SplitProtocol/Update/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1868/SplitProtocol/Update/cr
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1862/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1862/SplitProtocol/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1862/SplitProtocol/Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1862/SplitProtocol/Sample/rr
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1862/SplitProtocol/Update/$entry
      -- CP-element group 225: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1862/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1850_branch_ack_0, ack => zeropad3D_CP_2152_elements(225)); -- 
    rr_11616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(225), ack => type_cast_1868_inst_req_0); -- 
    cr_11621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(225), ack => type_cast_1868_inst_req_1); -- 
    rr_11639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(225), ack => type_cast_1862_inst_req_0); -- 
    cr_11644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(225), ack => type_cast_1862_inst_req_1); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	889 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1890_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1890_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1890_Sample/ra
      -- 
    ra_4948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1890_inst_ack_0, ack => zeropad3D_CP_2152_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	889 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	240 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1890_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1890_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1890_Update/ca
      -- 
    ca_4953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1890_inst_ack_1, ack => zeropad3D_CP_2152_elements(227)); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	889 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (5) 
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Sample/word_access_start/$exit
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Sample/word_access_start/word_0/$exit
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Sample/word_access_start/word_0/ra
      -- 
    ra_4970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1899_load_0_ack_0, ack => zeropad3D_CP_2152_elements(228)); -- 
    -- CP-element group 229:  transition  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	889 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	238 
    -- CP-element group 229:  members (12) 
      -- CP-element group 229: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Update/word_access_complete/$exit
      -- CP-element group 229: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Update/word_access_complete/word_0/$exit
      -- CP-element group 229: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Update/word_access_complete/word_0/ca
      -- CP-element group 229: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Update/LOAD_pad_1899_Merge/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Update/LOAD_pad_1899_Merge/$exit
      -- CP-element group 229: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Update/LOAD_pad_1899_Merge/merge_req
      -- CP-element group 229: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Update/LOAD_pad_1899_Merge/merge_ack
      -- CP-element group 229: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1969_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1969_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1969_Sample/rr
      -- 
    ca_4981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1899_load_0_ack_1, ack => zeropad3D_CP_2152_elements(229)); -- 
    rr_5141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(229), ack => type_cast_1969_inst_req_0); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	889 
    -- CP-element group 230: successors 
    -- CP-element group 230:  members (5) 
      -- CP-element group 230: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_sample_completed_
      -- CP-element group 230: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Sample/word_access_start/$exit
      -- CP-element group 230: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Sample/word_access_start/word_0/$exit
      -- CP-element group 230: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Sample/word_access_start/word_0/ra
      -- 
    ra_5003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_1902_load_0_ack_0, ack => zeropad3D_CP_2152_elements(230)); -- 
    -- CP-element group 231:  transition  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	889 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	236 
    -- CP-element group 231:  members (12) 
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Update/word_access_complete/$exit
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Update/word_access_complete/word_0/$exit
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Update/word_access_complete/word_0/ca
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Update/LOAD_depth_high_1902_Merge/$entry
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Update/LOAD_depth_high_1902_Merge/$exit
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Update/LOAD_depth_high_1902_Merge/merge_req
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Update/LOAD_depth_high_1902_Merge/merge_ack
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1930_sample_start_
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1930_Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1930_Sample/rr
      -- 
    ca_5014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_1902_load_0_ack_1, ack => zeropad3D_CP_2152_elements(231)); -- 
    rr_5127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(231), ack => type_cast_1930_inst_req_0); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	889 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (5) 
      -- CP-element group 232: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Sample/word_access_start/$exit
      -- CP-element group 232: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Sample/word_access_start/word_0/$exit
      -- CP-element group 232: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Sample/word_access_start/word_0/ra
      -- 
    ra_5053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1914_load_0_ack_0, ack => zeropad3D_CP_2152_elements(232)); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	889 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	240 
    -- CP-element group 233:  members (9) 
      -- CP-element group 233: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Update/word_access_complete/$exit
      -- CP-element group 233: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Update/word_access_complete/word_0/$exit
      -- CP-element group 233: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Update/word_access_complete/word_0/ca
      -- CP-element group 233: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Update/ptr_deref_1914_Merge/$entry
      -- CP-element group 233: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Update/ptr_deref_1914_Merge/$exit
      -- CP-element group 233: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Update/ptr_deref_1914_Merge/merge_req
      -- CP-element group 233: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Update/ptr_deref_1914_Merge/merge_ack
      -- 
    ca_5064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1914_load_0_ack_1, ack => zeropad3D_CP_2152_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	889 
    -- CP-element group 234: successors 
    -- CP-element group 234:  members (5) 
      -- CP-element group 234: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_sample_completed_
      -- CP-element group 234: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Sample/word_access_start/$exit
      -- CP-element group 234: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Sample/word_access_start/word_0/$exit
      -- CP-element group 234: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Sample/word_access_start/word_0/ra
      -- 
    ra_5103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1926_load_0_ack_0, ack => zeropad3D_CP_2152_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	889 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	240 
    -- CP-element group 235:  members (9) 
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_update_completed_
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Update/word_access_complete/$exit
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Update/word_access_complete/word_0/$exit
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Update/word_access_complete/word_0/ca
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Update/ptr_deref_1926_Merge/$entry
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Update/ptr_deref_1926_Merge/$exit
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Update/ptr_deref_1926_Merge/merge_req
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Update/ptr_deref_1926_Merge/merge_ack
      -- 
    ca_5114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1926_load_0_ack_1, ack => zeropad3D_CP_2152_elements(235)); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	231 
    -- CP-element group 236: successors 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1930_sample_completed_
      -- CP-element group 236: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1930_Sample/$exit
      -- CP-element group 236: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1930_Sample/ra
      -- 
    ra_5128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1930_inst_ack_0, ack => zeropad3D_CP_2152_elements(236)); -- 
    -- CP-element group 237:  transition  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	889 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	240 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1930_update_completed_
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1930_Update/$exit
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1930_Update/ca
      -- 
    ca_5133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1930_inst_ack_1, ack => zeropad3D_CP_2152_elements(237)); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	229 
    -- CP-element group 238: successors 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1969_sample_completed_
      -- CP-element group 238: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1969_Sample/$exit
      -- CP-element group 238: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1969_Sample/ra
      -- 
    ra_5142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1969_inst_ack_0, ack => zeropad3D_CP_2152_elements(238)); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	889 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1969_update_completed_
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1969_Update/$exit
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1969_Update/ca
      -- 
    ca_5147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1969_inst_ack_1, ack => zeropad3D_CP_2152_elements(239)); -- 
    -- CP-element group 240:  join  fork  transition  place  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	227 
    -- CP-element group 240: 	233 
    -- CP-element group 240: 	235 
    -- CP-element group 240: 	237 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	900 
    -- CP-element group 240: 	901 
    -- CP-element group 240: 	902 
    -- CP-element group 240: 	903 
    -- CP-element group 240:  members (16) 
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460
      -- CP-element group 240: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011__exit__
      -- CP-element group 240: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/$exit
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/$entry
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2027/$entry
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/$entry
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2014/$entry
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/$entry
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/$entry
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/$entry
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2024/$entry
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2024/SplitProtocol/$entry
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2024/SplitProtocol/Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2024/SplitProtocol/Sample/rr
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2024/SplitProtocol/Update/$entry
      -- CP-element group 240: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2024/SplitProtocol/Update/cr
      -- 
    rr_11887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(240), ack => type_cast_2024_inst_req_0); -- 
    cr_11892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(240), ack => type_cast_2024_inst_req_1); -- 
    zeropad3D_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(227) & zeropad3D_CP_2152_elements(233) & zeropad3D_CP_2152_elements(235) & zeropad3D_CP_2152_elements(237) & zeropad3D_CP_2152_elements(239);
      gj_zeropad3D_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	910 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/type_cast_2038_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/type_cast_2038_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/type_cast_2038_Sample/ra
      -- 
    ra_5159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2038_inst_ack_0, ack => zeropad3D_CP_2152_elements(241)); -- 
    -- CP-element group 242:  branch  transition  place  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	910 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (13) 
      -- CP-element group 242: 	 branch_block_stmt_714/if_stmt_2047__entry__
      -- CP-element group 242: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046__exit__
      -- CP-element group 242: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/$exit
      -- CP-element group 242: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/type_cast_2038_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/type_cast_2038_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/type_cast_2038_Update/ca
      -- CP-element group 242: 	 branch_block_stmt_714/if_stmt_2047_dead_link/$entry
      -- CP-element group 242: 	 branch_block_stmt_714/if_stmt_2047_eval_test/$entry
      -- CP-element group 242: 	 branch_block_stmt_714/if_stmt_2047_eval_test/$exit
      -- CP-element group 242: 	 branch_block_stmt_714/if_stmt_2047_eval_test/branch_req
      -- CP-element group 242: 	 branch_block_stmt_714/R_cmp465_2048_place
      -- CP-element group 242: 	 branch_block_stmt_714/if_stmt_2047_if_link/$entry
      -- CP-element group 242: 	 branch_block_stmt_714/if_stmt_2047_else_link/$entry
      -- 
    ca_5164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2038_inst_ack_1, ack => zeropad3D_CP_2152_elements(242)); -- 
    branch_req_5172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(242), ack => if_stmt_2047_branch_req_0); -- 
    -- CP-element group 243:  transition  place  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	911 
    -- CP-element group 243:  members (5) 
      -- CP-element group 243: 	 branch_block_stmt_714/if_stmt_2047_if_link/$exit
      -- CP-element group 243: 	 branch_block_stmt_714/if_stmt_2047_if_link/if_choice_transition
      -- CP-element group 243: 	 branch_block_stmt_714/whilex_xbody460_ifx_xthen496
      -- CP-element group 243: 	 branch_block_stmt_714/whilex_xbody460_ifx_xthen496_PhiReq/$entry
      -- CP-element group 243: 	 branch_block_stmt_714/whilex_xbody460_ifx_xthen496_PhiReq/$exit
      -- 
    if_choice_transition_5177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2047_branch_ack_1, ack => zeropad3D_CP_2152_elements(243)); -- 
    -- CP-element group 244:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244: 	246 
    -- CP-element group 244: 	248 
    -- CP-element group 244:  members (27) 
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078__entry__
      -- CP-element group 244: 	 branch_block_stmt_714/merge_stmt_2053__exit__
      -- CP-element group 244: 	 branch_block_stmt_714/if_stmt_2047_else_link/$exit
      -- CP-element group 244: 	 branch_block_stmt_714/if_stmt_2047_else_link/else_choice_transition
      -- CP-element group 244: 	 branch_block_stmt_714/whilex_xbody460_lorx_xlhsx_xfalse467
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/$entry
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_update_start_
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_word_address_calculated
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_root_address_calculated
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Sample/word_access_start/$entry
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Sample/word_access_start/word_0/$entry
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Sample/word_access_start/word_0/rr
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Update/$entry
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Update/word_access_complete/$entry
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Update/word_access_complete/word_0/$entry
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Update/word_access_complete/word_0/cr
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/type_cast_2059_update_start_
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/type_cast_2059_Update/$entry
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/type_cast_2059_Update/cr
      -- CP-element group 244: 	 branch_block_stmt_714/whilex_xbody460_lorx_xlhsx_xfalse467_PhiReq/$entry
      -- CP-element group 244: 	 branch_block_stmt_714/whilex_xbody460_lorx_xlhsx_xfalse467_PhiReq/$exit
      -- CP-element group 244: 	 branch_block_stmt_714/merge_stmt_2053_PhiReqMerge
      -- CP-element group 244: 	 branch_block_stmt_714/merge_stmt_2053_PhiAck/$entry
      -- CP-element group 244: 	 branch_block_stmt_714/merge_stmt_2053_PhiAck/$exit
      -- CP-element group 244: 	 branch_block_stmt_714/merge_stmt_2053_PhiAck/dummy
      -- 
    else_choice_transition_5181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2047_branch_ack_0, ack => zeropad3D_CP_2152_elements(244)); -- 
    rr_5202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(244), ack => LOAD_row_high_2055_load_0_req_0); -- 
    cr_5213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(244), ack => LOAD_row_high_2055_load_0_req_1); -- 
    cr_5232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(244), ack => type_cast_2059_inst_req_1); -- 
    -- CP-element group 245:  transition  input  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245:  members (5) 
      -- CP-element group 245: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Sample/word_access_start/$exit
      -- CP-element group 245: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Sample/word_access_start/word_0/$exit
      -- CP-element group 245: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Sample/word_access_start/word_0/ra
      -- 
    ra_5203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2055_load_0_ack_0, ack => zeropad3D_CP_2152_elements(245)); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	244 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (12) 
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Update/word_access_complete/$exit
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Update/word_access_complete/word_0/$exit
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Update/word_access_complete/word_0/ca
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Update/LOAD_row_high_2055_Merge/$entry
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Update/LOAD_row_high_2055_Merge/$exit
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Update/LOAD_row_high_2055_Merge/merge_req
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/LOAD_row_high_2055_Update/LOAD_row_high_2055_Merge/merge_ack
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/type_cast_2059_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/type_cast_2059_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/type_cast_2059_Sample/rr
      -- 
    ca_5214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2055_load_0_ack_1, ack => zeropad3D_CP_2152_elements(246)); -- 
    rr_5227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(246), ack => type_cast_2059_inst_req_0); -- 
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/type_cast_2059_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/type_cast_2059_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/type_cast_2059_Sample/ra
      -- 
    ra_5228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2059_inst_ack_0, ack => zeropad3D_CP_2152_elements(247)); -- 
    -- CP-element group 248:  branch  transition  place  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	244 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248: 	250 
    -- CP-element group 248:  members (13) 
      -- CP-element group 248: 	 branch_block_stmt_714/if_stmt_2079__entry__
      -- CP-element group 248: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078__exit__
      -- CP-element group 248: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/$exit
      -- CP-element group 248: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/type_cast_2059_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/type_cast_2059_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_714/assign_stmt_2056_to_assign_stmt_2078/type_cast_2059_Update/ca
      -- CP-element group 248: 	 branch_block_stmt_714/if_stmt_2079_dead_link/$entry
      -- CP-element group 248: 	 branch_block_stmt_714/if_stmt_2079_eval_test/$entry
      -- CP-element group 248: 	 branch_block_stmt_714/if_stmt_2079_eval_test/$exit
      -- CP-element group 248: 	 branch_block_stmt_714/if_stmt_2079_eval_test/branch_req
      -- CP-element group 248: 	 branch_block_stmt_714/R_cmp476_2080_place
      -- CP-element group 248: 	 branch_block_stmt_714/if_stmt_2079_if_link/$entry
      -- CP-element group 248: 	 branch_block_stmt_714/if_stmt_2079_else_link/$entry
      -- 
    ca_5233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2059_inst_ack_1, ack => zeropad3D_CP_2152_elements(248)); -- 
    branch_req_5241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(248), ack => if_stmt_2079_branch_req_0); -- 
    -- CP-element group 249:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: 	252 
    -- CP-element group 249:  members (18) 
      -- CP-element group 249: 	 branch_block_stmt_714/merge_stmt_2085__exit__
      -- CP-element group 249: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097__entry__
      -- CP-element group 249: 	 branch_block_stmt_714/if_stmt_2079_if_link/$exit
      -- CP-element group 249: 	 branch_block_stmt_714/if_stmt_2079_if_link/if_choice_transition
      -- CP-element group 249: 	 branch_block_stmt_714/lorx_xlhsx_xfalse467_lorx_xlhsx_xfalse478
      -- CP-element group 249: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/$entry
      -- CP-element group 249: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/type_cast_2089_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/type_cast_2089_update_start_
      -- CP-element group 249: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/type_cast_2089_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/type_cast_2089_Sample/rr
      -- CP-element group 249: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/type_cast_2089_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/type_cast_2089_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_714/lorx_xlhsx_xfalse467_lorx_xlhsx_xfalse478_PhiReq/$entry
      -- CP-element group 249: 	 branch_block_stmt_714/lorx_xlhsx_xfalse467_lorx_xlhsx_xfalse478_PhiReq/$exit
      -- CP-element group 249: 	 branch_block_stmt_714/merge_stmt_2085_PhiReqMerge
      -- CP-element group 249: 	 branch_block_stmt_714/merge_stmt_2085_PhiAck/$entry
      -- CP-element group 249: 	 branch_block_stmt_714/merge_stmt_2085_PhiAck/$exit
      -- CP-element group 249: 	 branch_block_stmt_714/merge_stmt_2085_PhiAck/dummy
      -- 
    if_choice_transition_5246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2079_branch_ack_1, ack => zeropad3D_CP_2152_elements(249)); -- 
    rr_5263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(249), ack => type_cast_2089_inst_req_0); -- 
    cr_5268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(249), ack => type_cast_2089_inst_req_1); -- 
    -- CP-element group 250:  transition  place  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	248 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	911 
    -- CP-element group 250:  members (5) 
      -- CP-element group 250: 	 branch_block_stmt_714/if_stmt_2079_else_link/$exit
      -- CP-element group 250: 	 branch_block_stmt_714/if_stmt_2079_else_link/else_choice_transition
      -- CP-element group 250: 	 branch_block_stmt_714/lorx_xlhsx_xfalse467_ifx_xthen496
      -- CP-element group 250: 	 branch_block_stmt_714/lorx_xlhsx_xfalse467_ifx_xthen496_PhiReq/$entry
      -- CP-element group 250: 	 branch_block_stmt_714/lorx_xlhsx_xfalse467_ifx_xthen496_PhiReq/$exit
      -- 
    else_choice_transition_5250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2079_branch_ack_0, ack => zeropad3D_CP_2152_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/type_cast_2089_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/type_cast_2089_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/type_cast_2089_Sample/ra
      -- 
    ra_5264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2089_inst_ack_0, ack => zeropad3D_CP_2152_elements(251)); -- 
    -- CP-element group 252:  branch  transition  place  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	249 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (13) 
      -- CP-element group 252: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097__exit__
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2098__entry__
      -- CP-element group 252: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/$exit
      -- CP-element group 252: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/type_cast_2089_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/type_cast_2089_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_714/assign_stmt_2090_to_assign_stmt_2097/type_cast_2089_Update/ca
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2098_dead_link/$entry
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2098_eval_test/$entry
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2098_eval_test/$exit
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2098_eval_test/branch_req
      -- CP-element group 252: 	 branch_block_stmt_714/R_cmp483_2099_place
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2098_if_link/$entry
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2098_else_link/$entry
      -- 
    ca_5269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2089_inst_ack_1, ack => zeropad3D_CP_2152_elements(252)); -- 
    branch_req_5277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(252), ack => if_stmt_2098_branch_req_0); -- 
    -- CP-element group 253:  transition  place  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	911 
    -- CP-element group 253:  members (5) 
      -- CP-element group 253: 	 branch_block_stmt_714/if_stmt_2098_if_link/$exit
      -- CP-element group 253: 	 branch_block_stmt_714/if_stmt_2098_if_link/if_choice_transition
      -- CP-element group 253: 	 branch_block_stmt_714/lorx_xlhsx_xfalse478_ifx_xthen496
      -- CP-element group 253: 	 branch_block_stmt_714/lorx_xlhsx_xfalse478_ifx_xthen496_PhiReq/$entry
      -- CP-element group 253: 	 branch_block_stmt_714/lorx_xlhsx_xfalse478_ifx_xthen496_PhiReq/$exit
      -- 
    if_choice_transition_5282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2098_branch_ack_1, ack => zeropad3D_CP_2152_elements(253)); -- 
    -- CP-element group 254:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254: 	256 
    -- CP-element group 254: 	258 
    -- CP-element group 254:  members (27) 
      -- CP-element group 254: 	 branch_block_stmt_714/merge_stmt_2104__exit__
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129__entry__
      -- CP-element group 254: 	 branch_block_stmt_714/if_stmt_2098_else_link/$exit
      -- CP-element group 254: 	 branch_block_stmt_714/if_stmt_2098_else_link/else_choice_transition
      -- CP-element group 254: 	 branch_block_stmt_714/lorx_xlhsx_xfalse478_lorx_xlhsx_xfalse485
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_update_start_
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_word_address_calculated
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_root_address_calculated
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Sample/word_access_start/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Sample/word_access_start/word_0/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Sample/word_access_start/word_0/rr
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Update/word_access_complete/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Update/word_access_complete/word_0/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Update/word_access_complete/word_0/cr
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/type_cast_2110_update_start_
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/type_cast_2110_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/type_cast_2110_Update/cr
      -- CP-element group 254: 	 branch_block_stmt_714/lorx_xlhsx_xfalse478_lorx_xlhsx_xfalse485_PhiReq/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/lorx_xlhsx_xfalse478_lorx_xlhsx_xfalse485_PhiReq/$exit
      -- CP-element group 254: 	 branch_block_stmt_714/merge_stmt_2104_PhiReqMerge
      -- CP-element group 254: 	 branch_block_stmt_714/merge_stmt_2104_PhiAck/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/merge_stmt_2104_PhiAck/$exit
      -- CP-element group 254: 	 branch_block_stmt_714/merge_stmt_2104_PhiAck/dummy
      -- 
    else_choice_transition_5286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2098_branch_ack_0, ack => zeropad3D_CP_2152_elements(254)); -- 
    rr_5307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(254), ack => LOAD_col_high_2106_load_0_req_0); -- 
    cr_5318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(254), ack => LOAD_col_high_2106_load_0_req_1); -- 
    cr_5337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(254), ack => type_cast_2110_inst_req_1); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255:  members (5) 
      -- CP-element group 255: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Sample/word_access_start/$exit
      -- CP-element group 255: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Sample/word_access_start/word_0/$exit
      -- CP-element group 255: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Sample/word_access_start/word_0/ra
      -- 
    ra_5308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2106_load_0_ack_0, ack => zeropad3D_CP_2152_elements(255)); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (12) 
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Update/word_access_complete/$exit
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Update/word_access_complete/word_0/$exit
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Update/word_access_complete/word_0/ca
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Update/LOAD_col_high_2106_Merge/$entry
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Update/LOAD_col_high_2106_Merge/$exit
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Update/LOAD_col_high_2106_Merge/merge_req
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/LOAD_col_high_2106_Update/LOAD_col_high_2106_Merge/merge_ack
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/type_cast_2110_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/type_cast_2110_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/type_cast_2110_Sample/rr
      -- 
    ca_5319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2106_load_0_ack_1, ack => zeropad3D_CP_2152_elements(256)); -- 
    rr_5332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(256), ack => type_cast_2110_inst_req_0); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/type_cast_2110_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/type_cast_2110_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/type_cast_2110_Sample/ra
      -- 
    ra_5333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2110_inst_ack_0, ack => zeropad3D_CP_2152_elements(257)); -- 
    -- CP-element group 258:  branch  transition  place  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	254 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (13) 
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2130__entry__
      -- CP-element group 258: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129__exit__
      -- CP-element group 258: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/$exit
      -- CP-element group 258: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/type_cast_2110_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/type_cast_2110_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_714/assign_stmt_2107_to_assign_stmt_2129/type_cast_2110_Update/ca
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2130_dead_link/$entry
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2130_eval_test/$entry
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2130_eval_test/$exit
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2130_eval_test/branch_req
      -- CP-element group 258: 	 branch_block_stmt_714/R_cmp494_2131_place
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2130_if_link/$entry
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2130_else_link/$entry
      -- 
    ca_5338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2110_inst_ack_1, ack => zeropad3D_CP_2152_elements(258)); -- 
    branch_req_5346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(258), ack => if_stmt_2130_branch_req_0); -- 
    -- CP-element group 259:  fork  transition  place  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	275 
    -- CP-element group 259: 	276 
    -- CP-element group 259: 	278 
    -- CP-element group 259: 	280 
    -- CP-element group 259: 	282 
    -- CP-element group 259: 	284 
    -- CP-element group 259: 	286 
    -- CP-element group 259: 	288 
    -- CP-element group 259: 	290 
    -- CP-element group 259: 	293 
    -- CP-element group 259:  members (46) 
      -- CP-element group 259: 	 branch_block_stmt_714/merge_stmt_2194__exit__
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299__entry__
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_final_index_sum_regn_update_start
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2287_update_start_
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2262_update_start_
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2198_Update/cr
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2198_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2198_Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_update_start_
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Update/word_access_complete/word_0/cr
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Update/word_access_complete/word_0/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Update/word_access_complete/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2294_complete/req
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2294_complete/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Update/word_access_complete/word_0/cr
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Update/word_access_complete/word_0/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Update/word_access_complete/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2294_update_start_
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2198_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2198_update_start_
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2287_Update/cr
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2198_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2287_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_final_index_sum_regn_Update/req
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_final_index_sum_regn_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2269_update_start_
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_update_start_
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2269_complete/req
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2269_complete/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_final_index_sum_regn_update_start
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2262_Update/cr
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2262_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_final_index_sum_regn_Update/req
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_final_index_sum_regn_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/if_stmt_2130_if_link/$exit
      -- CP-element group 259: 	 branch_block_stmt_714/if_stmt_2130_if_link/if_choice_transition
      -- CP-element group 259: 	 branch_block_stmt_714/lorx_xlhsx_xfalse485_ifx_xelse517
      -- CP-element group 259: 	 branch_block_stmt_714/lorx_xlhsx_xfalse485_ifx_xelse517_PhiReq/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/lorx_xlhsx_xfalse485_ifx_xelse517_PhiReq/$exit
      -- CP-element group 259: 	 branch_block_stmt_714/merge_stmt_2194_PhiReqMerge
      -- CP-element group 259: 	 branch_block_stmt_714/merge_stmt_2194_PhiAck/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/merge_stmt_2194_PhiAck/$exit
      -- CP-element group 259: 	 branch_block_stmt_714/merge_stmt_2194_PhiAck/dummy
      -- 
    if_choice_transition_5351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2130_branch_ack_1, ack => zeropad3D_CP_2152_elements(259)); -- 
    cr_5514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(259), ack => type_cast_2198_inst_req_1); -- 
    rr_5509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(259), ack => type_cast_2198_inst_req_0); -- 
    cr_5734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(259), ack => ptr_deref_2297_store_0_req_1); -- 
    req_5684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(259), ack => addr_of_2294_final_reg_req_1); -- 
    cr_5619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(259), ack => ptr_deref_2273_load_0_req_1); -- 
    cr_5638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(259), ack => type_cast_2287_inst_req_1); -- 
    req_5669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(259), ack => array_obj_ref_2293_index_offset_req_1); -- 
    req_5574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(259), ack => addr_of_2269_final_reg_req_1); -- 
    cr_5528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(259), ack => type_cast_2262_inst_req_1); -- 
    req_5559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(259), ack => array_obj_ref_2268_index_offset_req_1); -- 
    -- CP-element group 260:  transition  place  input  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	911 
    -- CP-element group 260:  members (5) 
      -- CP-element group 260: 	 branch_block_stmt_714/if_stmt_2130_else_link/$exit
      -- CP-element group 260: 	 branch_block_stmt_714/if_stmt_2130_else_link/else_choice_transition
      -- CP-element group 260: 	 branch_block_stmt_714/lorx_xlhsx_xfalse485_ifx_xthen496
      -- CP-element group 260: 	 branch_block_stmt_714/lorx_xlhsx_xfalse485_ifx_xthen496_PhiReq/$entry
      -- CP-element group 260: 	 branch_block_stmt_714/lorx_xlhsx_xfalse485_ifx_xthen496_PhiReq/$exit
      -- 
    else_choice_transition_5355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2130_branch_ack_0, ack => zeropad3D_CP_2152_elements(260)); -- 
    -- CP-element group 261:  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	911 
    -- CP-element group 261: successors 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2140_sample_completed_
      -- CP-element group 261: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2140_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2140_Sample/ra
      -- 
    ra_5369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2140_inst_ack_0, ack => zeropad3D_CP_2152_elements(261)); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	911 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	265 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2140_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2140_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2140_Update/ca
      -- 
    ca_5374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2140_inst_ack_1, ack => zeropad3D_CP_2152_elements(262)); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	911 
    -- CP-element group 263: successors 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2145_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2145_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2145_Sample/ra
      -- 
    ra_5383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2145_inst_ack_0, ack => zeropad3D_CP_2152_elements(263)); -- 
    -- CP-element group 264:  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	911 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2145_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2145_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2145_Update/ca
      -- 
    ca_5388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2145_inst_ack_1, ack => zeropad3D_CP_2152_elements(264)); -- 
    -- CP-element group 265:  join  transition  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	262 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2179_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2179_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2179_Sample/rr
      -- 
    rr_5396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(265), ack => type_cast_2179_inst_req_0); -- 
    zeropad3D_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(262) & zeropad3D_CP_2152_elements(264);
      gj_zeropad3D_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2179_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2179_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2179_Sample/ra
      -- 
    ra_5397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2179_inst_ack_0, ack => zeropad3D_CP_2152_elements(266)); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	911 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (16) 
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2179_update_completed_
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2179_Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2179_Update/ca
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_index_resized_1
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_index_scaled_1
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_index_computed_1
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_index_resize_1/$entry
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_index_resize_1/$exit
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_index_resize_1/index_resize_req
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_index_resize_1/index_resize_ack
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_index_scale_1/$entry
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_index_scale_1/$exit
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_index_scale_1/scale_rename_req
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_index_scale_1/scale_rename_ack
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_final_index_sum_regn_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_final_index_sum_regn_Sample/req
      -- 
    ca_5402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2179_inst_ack_1, ack => zeropad3D_CP_2152_elements(267)); -- 
    req_5427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(267), ack => array_obj_ref_2185_index_offset_req_0); -- 
    -- CP-element group 268:  transition  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	274 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_final_index_sum_regn_sample_complete
      -- CP-element group 268: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_final_index_sum_regn_Sample/$exit
      -- CP-element group 268: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_final_index_sum_regn_Sample/ack
      -- 
    ack_5428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2185_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(268)); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	911 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (11) 
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/addr_of_2186_sample_start_
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_root_address_calculated
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_offset_calculated
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_final_index_sum_regn_Update/$exit
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_final_index_sum_regn_Update/ack
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_base_plus_offset/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_base_plus_offset/$exit
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_base_plus_offset/sum_rename_req
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_base_plus_offset/sum_rename_ack
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/addr_of_2186_request/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/addr_of_2186_request/req
      -- 
    ack_5433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2185_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(269)); -- 
    req_5442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(269), ack => addr_of_2186_final_reg_req_0); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/addr_of_2186_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/addr_of_2186_request/$exit
      -- CP-element group 270: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/addr_of_2186_request/ack
      -- 
    ack_5443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2186_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(270)); -- 
    -- CP-element group 271:  join  fork  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	911 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (28) 
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Sample/word_access_start/word_0/rr
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Sample/word_access_start/word_0/$entry
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Sample/word_access_start/$entry
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Sample/ptr_deref_2189_Split/split_ack
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Sample/ptr_deref_2189_Split/split_req
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/addr_of_2186_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/addr_of_2186_complete/$exit
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/addr_of_2186_complete/ack
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_sample_start_
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_base_address_calculated
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_word_address_calculated
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_root_address_calculated
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_base_address_resized
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_base_addr_resize/$entry
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_base_addr_resize/$exit
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_base_addr_resize/base_resize_req
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_base_addr_resize/base_resize_ack
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_base_plus_offset/$entry
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_base_plus_offset/$exit
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_base_plus_offset/sum_rename_req
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_base_plus_offset/sum_rename_ack
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_word_addrgen/$entry
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_word_addrgen/$exit
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_word_addrgen/root_register_req
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_word_addrgen/root_register_ack
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Sample/ptr_deref_2189_Split/$entry
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Sample/ptr_deref_2189_Split/$exit
      -- 
    ack_5448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2186_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(271)); -- 
    rr_5486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(271), ack => ptr_deref_2189_store_0_req_0); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (5) 
      -- CP-element group 272: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Sample/word_access_start/word_0/ra
      -- CP-element group 272: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Sample/word_access_start/word_0/$exit
      -- CP-element group 272: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Sample/word_access_start/$exit
      -- CP-element group 272: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Sample/$exit
      -- 
    ra_5487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2189_store_0_ack_0, ack => zeropad3D_CP_2152_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	911 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (5) 
      -- CP-element group 273: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Update/word_access_complete/word_0/$exit
      -- CP-element group 273: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Update/word_access_complete/word_0/ca
      -- CP-element group 273: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Update/word_access_complete/$exit
      -- CP-element group 273: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_update_completed_
      -- 
    ca_5498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2189_store_0_ack_1, ack => zeropad3D_CP_2152_elements(273)); -- 
    -- CP-element group 274:  join  transition  place  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: 	268 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	912 
    -- CP-element group 274:  members (5) 
      -- CP-element group 274: 	 branch_block_stmt_714/ifx_xthen496_ifx_xend565
      -- CP-element group 274: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192__exit__
      -- CP-element group 274: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/$exit
      -- CP-element group 274: 	 branch_block_stmt_714/ifx_xthen496_ifx_xend565_PhiReq/$entry
      -- CP-element group 274: 	 branch_block_stmt_714/ifx_xthen496_ifx_xend565_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(273) & zeropad3D_CP_2152_elements(268);
      gj_zeropad3D_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	259 
    -- CP-element group 275: successors 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2198_Sample/ra
      -- CP-element group 275: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2198_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2198_sample_completed_
      -- 
    ra_5510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2198_inst_ack_0, ack => zeropad3D_CP_2152_elements(275)); -- 
    -- CP-element group 276:  fork  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	259 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276: 	285 
    -- CP-element group 276:  members (9) 
      -- CP-element group 276: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2287_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2262_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2198_Update/ca
      -- CP-element group 276: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2198_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2198_update_completed_
      -- CP-element group 276: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2262_Sample/rr
      -- CP-element group 276: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2262_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2287_Sample/rr
      -- CP-element group 276: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2287_Sample/$entry
      -- 
    ca_5515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2198_inst_ack_1, ack => zeropad3D_CP_2152_elements(276)); -- 
    rr_5523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(276), ack => type_cast_2262_inst_req_0); -- 
    rr_5633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(276), ack => type_cast_2287_inst_req_0); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2262_sample_completed_
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2262_Sample/ra
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2262_Sample/$exit
      -- 
    ra_5524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2262_inst_ack_0, ack => zeropad3D_CP_2152_elements(277)); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	259 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (16) 
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2262_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_index_scale_1/scale_rename_ack
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_index_scale_1/scale_rename_req
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_index_scale_1/$exit
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_index_scale_1/$entry
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_index_resize_1/index_resize_ack
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_index_resize_1/index_resize_req
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_index_resize_1/$exit
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_index_resize_1/$entry
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_index_computed_1
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_index_scaled_1
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2262_Update/ca
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2262_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_index_resized_1
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_final_index_sum_regn_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_final_index_sum_regn_Sample/$entry
      -- 
    ca_5529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2262_inst_ack_1, ack => zeropad3D_CP_2152_elements(278)); -- 
    req_5554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(278), ack => array_obj_ref_2268_index_offset_req_0); -- 
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	294 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_final_index_sum_regn_sample_complete
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_final_index_sum_regn_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_final_index_sum_regn_Sample/$exit
      -- 
    ack_5555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2268_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(279)); -- 
    -- CP-element group 280:  transition  input  output  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	259 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (11) 
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_root_address_calculated
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2269_sample_start_
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2269_request/req
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2269_request/$entry
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_base_plus_offset/sum_rename_ack
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_base_plus_offset/sum_rename_req
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_base_plus_offset/$exit
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_base_plus_offset/$entry
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_final_index_sum_regn_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_final_index_sum_regn_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2268_offset_calculated
      -- 
    ack_5560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2268_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(280)); -- 
    req_5569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(280), ack => addr_of_2269_final_reg_req_0); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2269_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2269_request/ack
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2269_request/$exit
      -- 
    ack_5570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2269_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(281)); -- 
    -- CP-element group 282:  join  fork  transition  input  output  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	259 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (24) 
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Sample/word_access_start/word_0/rr
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Sample/word_access_start/word_0/$entry
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Sample/word_access_start/$entry
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Sample/$entry
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_word_addrgen/root_register_ack
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_word_addrgen/root_register_req
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_word_addrgen/$exit
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_word_addrgen/$entry
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_base_plus_offset/sum_rename_ack
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_base_plus_offset/sum_rename_req
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_base_plus_offset/$exit
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_base_plus_offset/$entry
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_base_addr_resize/base_resize_ack
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2269_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_base_addr_resize/base_resize_req
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_base_addr_resize/$exit
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_base_addr_resize/$entry
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_base_address_resized
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_root_address_calculated
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_word_address_calculated
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_base_address_calculated
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_sample_start_
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2269_complete/ack
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2269_complete/$exit
      -- 
    ack_5575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2269_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(282)); -- 
    rr_5608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(282), ack => ptr_deref_2273_load_0_req_0); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283:  members (5) 
      -- CP-element group 283: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Sample/word_access_start/word_0/ra
      -- CP-element group 283: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Sample/word_access_start/word_0/$exit
      -- CP-element group 283: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Sample/word_access_start/$exit
      -- CP-element group 283: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_sample_completed_
      -- 
    ra_5609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2273_load_0_ack_0, ack => zeropad3D_CP_2152_elements(283)); -- 
    -- CP-element group 284:  transition  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	259 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	291 
    -- CP-element group 284:  members (9) 
      -- CP-element group 284: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Update/ptr_deref_2273_Merge/merge_ack
      -- CP-element group 284: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Update/ptr_deref_2273_Merge/merge_req
      -- CP-element group 284: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Update/ptr_deref_2273_Merge/$exit
      -- CP-element group 284: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Update/ptr_deref_2273_Merge/$entry
      -- CP-element group 284: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Update/word_access_complete/word_0/ca
      -- CP-element group 284: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Update/word_access_complete/word_0/$exit
      -- CP-element group 284: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Update/word_access_complete/$exit
      -- CP-element group 284: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2273_update_completed_
      -- 
    ca_5620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2273_load_0_ack_1, ack => zeropad3D_CP_2152_elements(284)); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	276 
    -- CP-element group 285: successors 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2287_sample_completed_
      -- CP-element group 285: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2287_Sample/ra
      -- CP-element group 285: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2287_Sample/$exit
      -- 
    ra_5634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2287_inst_ack_0, ack => zeropad3D_CP_2152_elements(285)); -- 
    -- CP-element group 286:  transition  input  output  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	259 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (16) 
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_index_resized_1
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_index_scaled_1
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_index_computed_1
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2287_Update/ca
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2287_Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_final_index_sum_regn_Sample/req
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_final_index_sum_regn_Sample/$entry
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_index_scale_1/scale_rename_ack
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_index_scale_1/scale_rename_req
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_index_scale_1/$exit
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_index_scale_1/$entry
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_index_resize_1/index_resize_ack
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_index_resize_1/index_resize_req
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_index_resize_1/$exit
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/type_cast_2287_update_completed_
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_index_resize_1/$entry
      -- 
    ca_5639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2287_inst_ack_1, ack => zeropad3D_CP_2152_elements(286)); -- 
    req_5664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(286), ack => array_obj_ref_2293_index_offset_req_0); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	294 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_final_index_sum_regn_Sample/ack
      -- CP-element group 287: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_final_index_sum_regn_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_final_index_sum_regn_sample_complete
      -- 
    ack_5665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2293_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(287)); -- 
    -- CP-element group 288:  transition  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	259 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (11) 
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_offset_calculated
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_root_address_calculated
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2294_request/req
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2294_request/$entry
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_base_plus_offset/sum_rename_ack
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2294_sample_start_
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_base_plus_offset/sum_rename_req
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_base_plus_offset/$exit
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_base_plus_offset/$entry
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_final_index_sum_regn_Update/ack
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/array_obj_ref_2293_final_index_sum_regn_Update/$exit
      -- 
    ack_5670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2293_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(288)); -- 
    req_5679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(288), ack => addr_of_2294_final_reg_req_0); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2294_request/ack
      -- CP-element group 289: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2294_sample_completed_
      -- CP-element group 289: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2294_request/$exit
      -- 
    ack_5680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2294_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(289)); -- 
    -- CP-element group 290:  fork  transition  input  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	259 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (19) 
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_base_addr_resize/$entry
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_base_addr_resize/$exit
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_base_addr_resize/base_resize_req
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_base_addr_resize/base_resize_ack
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_base_address_resized
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_root_address_calculated
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_word_address_calculated
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_base_address_calculated
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2294_complete/ack
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2294_complete/$exit
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/addr_of_2294_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_word_addrgen/root_register_ack
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_word_addrgen/root_register_req
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_word_addrgen/$exit
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_word_addrgen/$entry
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_base_plus_offset/sum_rename_ack
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_base_plus_offset/sum_rename_req
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_base_plus_offset/$exit
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_base_plus_offset/$entry
      -- 
    ack_5685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2294_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(290)); -- 
    -- CP-element group 291:  join  transition  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	284 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (9) 
      -- CP-element group 291: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_sample_start_
      -- CP-element group 291: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Sample/word_access_start/word_0/rr
      -- CP-element group 291: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Sample/word_access_start/word_0/$entry
      -- CP-element group 291: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Sample/word_access_start/$entry
      -- CP-element group 291: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Sample/ptr_deref_2297_Split/split_ack
      -- CP-element group 291: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Sample/ptr_deref_2297_Split/split_req
      -- CP-element group 291: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Sample/ptr_deref_2297_Split/$exit
      -- CP-element group 291: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Sample/ptr_deref_2297_Split/$entry
      -- CP-element group 291: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Sample/$entry
      -- 
    rr_5723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(291), ack => ptr_deref_2297_store_0_req_0); -- 
    zeropad3D_cp_element_group_291: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_291"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(284) & zeropad3D_CP_2152_elements(290);
      gj_zeropad3D_cp_element_group_291 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(291), clk => clk, reset => reset); --
    end block;
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292:  members (5) 
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_sample_completed_
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Sample/word_access_start/word_0/ra
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Sample/word_access_start/word_0/$exit
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Sample/word_access_start/$exit
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Sample/$exit
      -- 
    ra_5724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2297_store_0_ack_0, ack => zeropad3D_CP_2152_elements(292)); -- 
    -- CP-element group 293:  transition  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	259 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (5) 
      -- CP-element group 293: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Update/word_access_complete/word_0/ca
      -- CP-element group 293: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_update_completed_
      -- CP-element group 293: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Update/word_access_complete/word_0/$exit
      -- CP-element group 293: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Update/word_access_complete/$exit
      -- CP-element group 293: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/ptr_deref_2297_Update/$exit
      -- 
    ca_5735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2297_store_0_ack_1, ack => zeropad3D_CP_2152_elements(293)); -- 
    -- CP-element group 294:  join  transition  place  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	279 
    -- CP-element group 294: 	287 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	912 
    -- CP-element group 294:  members (5) 
      -- CP-element group 294: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299__exit__
      -- CP-element group 294: 	 branch_block_stmt_714/ifx_xelse517_ifx_xend565
      -- CP-element group 294: 	 branch_block_stmt_714/assign_stmt_2199_to_assign_stmt_2299/$exit
      -- CP-element group 294: 	 branch_block_stmt_714/ifx_xelse517_ifx_xend565_PhiReq/$entry
      -- CP-element group 294: 	 branch_block_stmt_714/ifx_xelse517_ifx_xend565_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(279) & zeropad3D_CP_2152_elements(287) & zeropad3D_CP_2152_elements(293);
      gj_zeropad3D_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	912 
    -- CP-element group 295: successors 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/type_cast_2305_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/type_cast_2305_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/type_cast_2305_Sample/ra
      -- 
    ra_5747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2305_inst_ack_0, ack => zeropad3D_CP_2152_elements(295)); -- 
    -- CP-element group 296:  branch  transition  place  input  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	912 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296: 	298 
    -- CP-element group 296:  members (13) 
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319__exit__
      -- CP-element group 296: 	 branch_block_stmt_714/if_stmt_2320__entry__
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/type_cast_2305_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/$exit
      -- CP-element group 296: 	 branch_block_stmt_714/if_stmt_2320_else_link/$entry
      -- CP-element group 296: 	 branch_block_stmt_714/if_stmt_2320_if_link/$entry
      -- CP-element group 296: 	 branch_block_stmt_714/if_stmt_2320_eval_test/branch_req
      -- CP-element group 296: 	 branch_block_stmt_714/if_stmt_2320_eval_test/$exit
      -- CP-element group 296: 	 branch_block_stmt_714/if_stmt_2320_eval_test/$entry
      -- CP-element group 296: 	 branch_block_stmt_714/if_stmt_2320_dead_link/$entry
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/type_cast_2305_Update/ca
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/type_cast_2305_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_714/R_cmp573_2321_place
      -- 
    ca_5752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2305_inst_ack_1, ack => zeropad3D_CP_2152_elements(296)); -- 
    branch_req_5760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(296), ack => if_stmt_2320_branch_req_0); -- 
    -- CP-element group 297:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	921 
    -- CP-element group 297: 	922 
    -- CP-element group 297: 	924 
    -- CP-element group 297: 	925 
    -- CP-element group 297: 	927 
    -- CP-element group 297: 	928 
    -- CP-element group 297:  members (40) 
      -- CP-element group 297: 	 branch_block_stmt_714/assign_stmt_2332__exit__
      -- CP-element group 297: 	 branch_block_stmt_714/assign_stmt_2332__entry__
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617
      -- CP-element group 297: 	 branch_block_stmt_714/merge_stmt_2326__exit__
      -- CP-element group 297: 	 branch_block_stmt_714/assign_stmt_2332/$exit
      -- CP-element group 297: 	 branch_block_stmt_714/assign_stmt_2332/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/if_stmt_2320_if_link/if_choice_transition
      -- CP-element group 297: 	 branch_block_stmt_714/if_stmt_2320_if_link/$exit
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xend565_ifx_xthen575
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xend565_ifx_xthen575_PhiReq/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xend565_ifx_xthen575_PhiReq/$exit
      -- CP-element group 297: 	 branch_block_stmt_714/merge_stmt_2326_PhiReqMerge
      -- CP-element group 297: 	 branch_block_stmt_714/merge_stmt_2326_PhiAck/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/merge_stmt_2326_PhiAck/$exit
      -- CP-element group 297: 	 branch_block_stmt_714/merge_stmt_2326_PhiAck/dummy
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/type_cast_2423/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/type_cast_2423/SplitProtocol/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/type_cast_2423/SplitProtocol/Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/type_cast_2423/SplitProtocol/Sample/rr
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/type_cast_2423/SplitProtocol/Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/type_cast_2423/SplitProtocol/Update/cr
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2430/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2430/SplitProtocol/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2430/SplitProtocol/Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2430/SplitProtocol/Sample/rr
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2430/SplitProtocol/Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2430/SplitProtocol/Update/cr
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Sample/rr
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2320_branch_ack_1, ack => zeropad3D_CP_2152_elements(297)); -- 
    rr_12077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(297), ack => type_cast_2423_inst_req_0); -- 
    cr_12082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(297), ack => type_cast_2423_inst_req_1); -- 
    rr_12100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(297), ack => type_cast_2430_inst_req_0); -- 
    cr_12105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(297), ack => type_cast_2430_inst_req_1); -- 
    rr_12123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(297), ack => type_cast_2436_inst_req_0); -- 
    cr_12128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(297), ack => type_cast_2436_inst_req_1); -- 
    -- CP-element group 298:  fork  transition  place  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	296 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298: 	300 
    -- CP-element group 298: 	301 
    -- CP-element group 298: 	302 
    -- CP-element group 298: 	304 
    -- CP-element group 298: 	307 
    -- CP-element group 298: 	309 
    -- CP-element group 298: 	310 
    -- CP-element group 298: 	311 
    -- CP-element group 298: 	313 
    -- CP-element group 298:  members (54) 
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412__entry__
      -- CP-element group 298: 	 branch_block_stmt_714/merge_stmt_2334__exit__
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_update_start_
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2344_Sample/rr
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2344_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Update/word_access_complete/word_0/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Sample/word_access_start/word_0/rr
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2344_update_start_
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2344_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Sample/word_access_start/word_0/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/if_stmt_2320_else_link/else_choice_transition
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Sample/word_access_start/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/ifx_xend565_ifx_xelse580
      -- CP-element group 298: 	 branch_block_stmt_714/if_stmt_2320_else_link/$exit
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_root_address_calculated
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Update/word_access_complete/word_0/cr
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_word_address_calculated
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2344_Update/cr
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Update/word_access_complete/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2344_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2351_update_start_
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2351_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2351_Update/cr
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2371_update_start_
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2371_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2371_Update/cr
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2388_update_start_
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2388_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2388_Update/cr
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_update_start_
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_word_address_calculated
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_root_address_calculated
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Sample/word_access_start/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Sample/word_access_start/word_0/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Sample/word_access_start/word_0/rr
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Update/word_access_complete/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Update/word_access_complete/word_0/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Update/word_access_complete/word_0/cr
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2395_update_start_
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2395_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2395_Update/cr
      -- CP-element group 298: 	 branch_block_stmt_714/ifx_xend565_ifx_xelse580_PhiReq/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/ifx_xend565_ifx_xelse580_PhiReq/$exit
      -- CP-element group 298: 	 branch_block_stmt_714/merge_stmt_2334_PhiReqMerge
      -- CP-element group 298: 	 branch_block_stmt_714/merge_stmt_2334_PhiAck/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/merge_stmt_2334_PhiAck/$exit
      -- CP-element group 298: 	 branch_block_stmt_714/merge_stmt_2334_PhiAck/dummy
      -- 
    else_choice_transition_5769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2320_branch_ack_0, ack => zeropad3D_CP_2152_elements(298)); -- 
    rr_5785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(298), ack => type_cast_2344_inst_req_0); -- 
    rr_5807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(298), ack => LOAD_col_high_2347_load_0_req_0); -- 
    cr_5818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(298), ack => LOAD_col_high_2347_load_0_req_1); -- 
    cr_5790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(298), ack => type_cast_2344_inst_req_1); -- 
    cr_5837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(298), ack => type_cast_2351_inst_req_1); -- 
    cr_5851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(298), ack => type_cast_2371_inst_req_1); -- 
    cr_5865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(298), ack => type_cast_2388_inst_req_1); -- 
    rr_5882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(298), ack => LOAD_row_high_2391_load_0_req_0); -- 
    cr_5893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(298), ack => LOAD_row_high_2391_load_0_req_1); -- 
    cr_5912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(298), ack => type_cast_2395_inst_req_1); -- 
    -- CP-element group 299:  transition  input  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2344_Sample/ra
      -- CP-element group 299: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2344_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2344_sample_completed_
      -- 
    ra_5786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2344_inst_ack_0, ack => zeropad3D_CP_2152_elements(299)); -- 
    -- CP-element group 300:  transition  input  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	305 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2344_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2344_Update/ca
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2344_Update/$exit
      -- 
    ca_5791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2344_inst_ack_1, ack => zeropad3D_CP_2152_elements(300)); -- 
    -- CP-element group 301:  transition  input  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	298 
    -- CP-element group 301: successors 
    -- CP-element group 301:  members (5) 
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Sample/word_access_start/word_0/ra
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Sample/word_access_start/word_0/$exit
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_sample_completed_
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Sample/word_access_start/$exit
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Sample/$exit
      -- 
    ra_5808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2347_load_0_ack_0, ack => zeropad3D_CP_2152_elements(301)); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	298 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (12) 
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Update/LOAD_col_high_2347_Merge/$exit
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Update/word_access_complete/word_0/$exit
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Update/word_access_complete/$exit
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Update/word_access_complete/word_0/ca
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_update_completed_
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Update/LOAD_col_high_2347_Merge/$entry
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Update/LOAD_col_high_2347_Merge/merge_req
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_col_high_2347_Update/LOAD_col_high_2347_Merge/merge_ack
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2351_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2351_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2351_Sample/rr
      -- 
    ca_5819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2347_load_0_ack_1, ack => zeropad3D_CP_2152_elements(302)); -- 
    rr_5832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(302), ack => type_cast_2351_inst_req_0); -- 
    -- CP-element group 303:  transition  input  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2351_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2351_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2351_Sample/ra
      -- 
    ra_5833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_0, ack => zeropad3D_CP_2152_elements(303)); -- 
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	298 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2351_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2351_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2351_Update/ca
      -- 
    ca_5838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_1, ack => zeropad3D_CP_2152_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	300 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2371_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2371_Sample/$entry
      -- CP-element group 305: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2371_Sample/rr
      -- 
    rr_5846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(305), ack => type_cast_2371_inst_req_0); -- 
    zeropad3D_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(300) & zeropad3D_CP_2152_elements(304);
      gj_zeropad3D_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2371_sample_completed_
      -- CP-element group 306: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2371_Sample/$exit
      -- CP-element group 306: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2371_Sample/ra
      -- 
    ra_5847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2371_inst_ack_0, ack => zeropad3D_CP_2152_elements(306)); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	298 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2371_update_completed_
      -- CP-element group 307: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2371_Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2371_Update/ca
      -- CP-element group 307: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2388_sample_start_
      -- CP-element group 307: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2388_Sample/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2388_Sample/rr
      -- 
    ca_5852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2371_inst_ack_1, ack => zeropad3D_CP_2152_elements(307)); -- 
    rr_5860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(307), ack => type_cast_2388_inst_req_0); -- 
    -- CP-element group 308:  transition  input  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2388_sample_completed_
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2388_Sample/$exit
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2388_Sample/ra
      -- 
    ra_5861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2388_inst_ack_0, ack => zeropad3D_CP_2152_elements(308)); -- 
    -- CP-element group 309:  transition  input  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	298 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	314 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2388_update_completed_
      -- CP-element group 309: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2388_Update/$exit
      -- CP-element group 309: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2388_Update/ca
      -- 
    ca_5866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2388_inst_ack_1, ack => zeropad3D_CP_2152_elements(309)); -- 
    -- CP-element group 310:  transition  input  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	298 
    -- CP-element group 310: successors 
    -- CP-element group 310:  members (5) 
      -- CP-element group 310: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_sample_completed_
      -- CP-element group 310: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Sample/$exit
      -- CP-element group 310: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Sample/word_access_start/$exit
      -- CP-element group 310: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Sample/word_access_start/word_0/$exit
      -- CP-element group 310: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Sample/word_access_start/word_0/ra
      -- 
    ra_5883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2391_load_0_ack_0, ack => zeropad3D_CP_2152_elements(310)); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	298 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (12) 
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_update_completed_
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Update/$exit
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Update/word_access_complete/$exit
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Update/word_access_complete/word_0/$exit
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Update/word_access_complete/word_0/ca
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Update/LOAD_row_high_2391_Merge/$entry
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Update/LOAD_row_high_2391_Merge/$exit
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Update/LOAD_row_high_2391_Merge/merge_req
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/LOAD_row_high_2391_Update/LOAD_row_high_2391_Merge/merge_ack
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2395_sample_start_
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2395_Sample/$entry
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2395_Sample/rr
      -- 
    ca_5894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2391_load_0_ack_1, ack => zeropad3D_CP_2152_elements(311)); -- 
    rr_5907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(311), ack => type_cast_2395_inst_req_0); -- 
    -- CP-element group 312:  transition  input  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2395_sample_completed_
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2395_Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2395_Sample/ra
      -- 
    ra_5908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2395_inst_ack_0, ack => zeropad3D_CP_2152_elements(312)); -- 
    -- CP-element group 313:  transition  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	298 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2395_update_completed_
      -- CP-element group 313: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2395_Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/type_cast_2395_Update/ca
      -- 
    ca_5913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2395_inst_ack_1, ack => zeropad3D_CP_2152_elements(313)); -- 
    -- CP-element group 314:  branch  join  transition  place  output  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	309 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314: 	316 
    -- CP-element group 314:  members (10) 
      -- CP-element group 314: 	 branch_block_stmt_714/if_stmt_2413__entry__
      -- CP-element group 314: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412__exit__
      -- CP-element group 314: 	 branch_block_stmt_714/assign_stmt_2340_to_assign_stmt_2412/$exit
      -- CP-element group 314: 	 branch_block_stmt_714/R_cmp608_2414_place
      -- CP-element group 314: 	 branch_block_stmt_714/if_stmt_2413_dead_link/$entry
      -- CP-element group 314: 	 branch_block_stmt_714/if_stmt_2413_eval_test/$entry
      -- CP-element group 314: 	 branch_block_stmt_714/if_stmt_2413_eval_test/$exit
      -- CP-element group 314: 	 branch_block_stmt_714/if_stmt_2413_eval_test/branch_req
      -- CP-element group 314: 	 branch_block_stmt_714/if_stmt_2413_if_link/$entry
      -- CP-element group 314: 	 branch_block_stmt_714/if_stmt_2413_else_link/$entry
      -- 
    branch_req_5921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(314), ack => if_stmt_2413_branch_req_0); -- 
    zeropad3D_cp_element_group_314: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_314"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(309) & zeropad3D_CP_2152_elements(313);
      gj_zeropad3D_cp_element_group_314 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(314), clk => clk, reset => reset); --
    end block;
    -- CP-element group 315:  fork  transition  place  input  output  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	936 
    -- CP-element group 315: 	937 
    -- CP-element group 315: 	939 
    -- CP-element group 315: 	940 
    -- CP-element group 315: 	942 
    -- CP-element group 315: 	943 
    -- CP-element group 315:  members (28) 
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618
      -- CP-element group 315: 	 branch_block_stmt_714/if_stmt_2413_if_link/$exit
      -- CP-element group 315: 	 branch_block_stmt_714/if_stmt_2413_if_link/if_choice_transition
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/type_cast_2445/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/type_cast_2445/SplitProtocol/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/type_cast_2445/SplitProtocol/Sample/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/type_cast_2445/SplitProtocol/Sample/rr
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/type_cast_2445/SplitProtocol/Update/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/type_cast_2445/SplitProtocol/Update/cr
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Sample/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Sample/rr
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Update/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Update/cr
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/type_cast_2453/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/type_cast_2453/SplitProtocol/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/type_cast_2453/SplitProtocol/Sample/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/type_cast_2453/SplitProtocol/Sample/rr
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/type_cast_2453/SplitProtocol/Update/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/type_cast_2453/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2413_branch_ack_1, ack => zeropad3D_CP_2152_elements(315)); -- 
    rr_12156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(315), ack => type_cast_2445_inst_req_0); -- 
    cr_12161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(315), ack => type_cast_2445_inst_req_1); -- 
    rr_12179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(315), ack => type_cast_2449_inst_req_0); -- 
    cr_12184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(315), ack => type_cast_2449_inst_req_1); -- 
    rr_12202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(315), ack => type_cast_2453_inst_req_0); -- 
    cr_12207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(315), ack => type_cast_2453_inst_req_1); -- 
    -- CP-element group 316:  fork  transition  place  input  output  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	314 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	913 
    -- CP-element group 316: 	914 
    -- CP-element group 316: 	915 
    -- CP-element group 316: 	917 
    -- CP-element group 316: 	918 
    -- CP-element group 316:  members (22) 
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617
      -- CP-element group 316: 	 branch_block_stmt_714/if_stmt_2413_else_link/$exit
      -- CP-element group 316: 	 branch_block_stmt_714/if_stmt_2413_else_link/else_choice_transition
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2420/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2432/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2432/SplitProtocol/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2432/SplitProtocol/Sample/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2432/SplitProtocol/Sample/rr
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2432/SplitProtocol/Update/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2432/SplitProtocol/Update/cr
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Sample/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Sample/rr
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Update/$entry
      -- CP-element group 316: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2413_branch_ack_0, ack => zeropad3D_CP_2152_elements(316)); -- 
    rr_12028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(316), ack => type_cast_2432_inst_req_0); -- 
    cr_12033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(316), ack => type_cast_2432_inst_req_1); -- 
    rr_12051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(316), ack => type_cast_2438_inst_req_0); -- 
    cr_12056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(316), ack => type_cast_2438_inst_req_1); -- 
    -- CP-element group 317:  transition  input  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	949 
    -- CP-element group 317: successors 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2457_sample_completed_
      -- CP-element group 317: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2457_Sample/$exit
      -- CP-element group 317: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2457_Sample/ra
      -- 
    ra_5944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2457_inst_ack_0, ack => zeropad3D_CP_2152_elements(317)); -- 
    -- CP-element group 318:  transition  input  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	949 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	333 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2457_update_completed_
      -- CP-element group 318: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2457_Update/$exit
      -- CP-element group 318: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2457_Update/ca
      -- 
    ca_5949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2457_inst_ack_1, ack => zeropad3D_CP_2152_elements(318)); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	949 
    -- CP-element group 319: successors 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2467_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2467_Sample/$exit
      -- CP-element group 319: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2467_Sample/ra
      -- 
    ra_5958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2467_inst_ack_0, ack => zeropad3D_CP_2152_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	949 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	333 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2467_update_completed_
      -- CP-element group 320: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2467_Update/$exit
      -- CP-element group 320: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2467_Update/ca
      -- 
    ca_5963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2467_inst_ack_1, ack => zeropad3D_CP_2152_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	949 
    -- CP-element group 321: successors 
    -- CP-element group 321:  members (5) 
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_sample_completed_
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Sample/$exit
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Sample/word_access_start/$exit
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Sample/word_access_start/word_0/$exit
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Sample/word_access_start/word_0/ra
      -- 
    ra_5980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2476_load_0_ack_0, ack => zeropad3D_CP_2152_elements(321)); -- 
    -- CP-element group 322:  transition  input  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	949 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	331 
    -- CP-element group 322:  members (12) 
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_update_completed_
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Update/$exit
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Update/word_access_complete/$exit
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Update/word_access_complete/word_0/$exit
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Update/word_access_complete/word_0/ca
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Update/LOAD_pad_2476_Merge/$entry
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Update/LOAD_pad_2476_Merge/$exit
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Update/LOAD_pad_2476_Merge/merge_req
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Update/LOAD_pad_2476_Merge/merge_ack
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2546_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2546_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2546_Sample/rr
      -- 
    ca_5991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2476_load_0_ack_1, ack => zeropad3D_CP_2152_elements(322)); -- 
    rr_6151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(322), ack => type_cast_2546_inst_req_0); -- 
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	949 
    -- CP-element group 323: successors 
    -- CP-element group 323:  members (5) 
      -- CP-element group 323: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Sample/word_access_start/$exit
      -- CP-element group 323: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Sample/word_access_start/word_0/$exit
      -- CP-element group 323: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Sample/word_access_start/word_0/ra
      -- 
    ra_6013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_2479_load_0_ack_0, ack => zeropad3D_CP_2152_elements(323)); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	949 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	329 
    -- CP-element group 324:  members (12) 
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Update/word_access_complete/$exit
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Update/word_access_complete/word_0/$exit
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Update/word_access_complete/word_0/ca
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Update/LOAD_depth_high_2479_Merge/$entry
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Update/LOAD_depth_high_2479_Merge/$exit
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Update/LOAD_depth_high_2479_Merge/merge_req
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Update/LOAD_depth_high_2479_Merge/merge_ack
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2507_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2507_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2507_Sample/rr
      -- 
    ca_6024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_2479_load_0_ack_1, ack => zeropad3D_CP_2152_elements(324)); -- 
    rr_6137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(324), ack => type_cast_2507_inst_req_0); -- 
    -- CP-element group 325:  transition  input  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	949 
    -- CP-element group 325: successors 
    -- CP-element group 325:  members (5) 
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Sample/word_access_start/$exit
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Sample/word_access_start/word_0/$exit
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Sample/word_access_start/word_0/ra
      -- 
    ra_6063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2491_load_0_ack_0, ack => zeropad3D_CP_2152_elements(325)); -- 
    -- CP-element group 326:  transition  input  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	949 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	333 
    -- CP-element group 326:  members (9) 
      -- CP-element group 326: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Update/word_access_complete/$exit
      -- CP-element group 326: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Update/word_access_complete/word_0/$exit
      -- CP-element group 326: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Update/word_access_complete/word_0/ca
      -- CP-element group 326: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Update/ptr_deref_2491_Merge/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Update/ptr_deref_2491_Merge/$exit
      -- CP-element group 326: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Update/ptr_deref_2491_Merge/merge_req
      -- CP-element group 326: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Update/ptr_deref_2491_Merge/merge_ack
      -- 
    ca_6074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2491_load_0_ack_1, ack => zeropad3D_CP_2152_elements(326)); -- 
    -- CP-element group 327:  transition  input  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	949 
    -- CP-element group 327: successors 
    -- CP-element group 327:  members (5) 
      -- CP-element group 327: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Sample/word_access_start/$exit
      -- CP-element group 327: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Sample/word_access_start/word_0/$exit
      -- CP-element group 327: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Sample/word_access_start/word_0/ra
      -- 
    ra_6113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2503_load_0_ack_0, ack => zeropad3D_CP_2152_elements(327)); -- 
    -- CP-element group 328:  transition  input  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	949 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	333 
    -- CP-element group 328:  members (9) 
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Update/word_access_complete/$exit
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Update/word_access_complete/word_0/$exit
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Update/word_access_complete/word_0/ca
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Update/ptr_deref_2503_Merge/$entry
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Update/ptr_deref_2503_Merge/$exit
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Update/ptr_deref_2503_Merge/merge_req
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Update/ptr_deref_2503_Merge/merge_ack
      -- 
    ca_6124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2503_load_0_ack_1, ack => zeropad3D_CP_2152_elements(328)); -- 
    -- CP-element group 329:  transition  input  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	324 
    -- CP-element group 329: successors 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2507_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2507_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2507_Sample/ra
      -- 
    ra_6138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2507_inst_ack_0, ack => zeropad3D_CP_2152_elements(329)); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	949 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	333 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2507_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2507_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2507_Update/ca
      -- 
    ca_6143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2507_inst_ack_1, ack => zeropad3D_CP_2152_elements(330)); -- 
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	322 
    -- CP-element group 331: successors 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2546_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2546_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2546_Sample/ra
      -- 
    ra_6152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2546_inst_ack_0, ack => zeropad3D_CP_2152_elements(331)); -- 
    -- CP-element group 332:  transition  input  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	949 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2546_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2546_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2546_Update/ca
      -- 
    ca_6157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2546_inst_ack_1, ack => zeropad3D_CP_2152_elements(332)); -- 
    -- CP-element group 333:  join  fork  transition  place  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	318 
    -- CP-element group 333: 	320 
    -- CP-element group 333: 	326 
    -- CP-element group 333: 	328 
    -- CP-element group 333: 	330 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	960 
    -- CP-element group 333: 	961 
    -- CP-element group 333: 	962 
    -- CP-element group 333: 	964 
    -- CP-element group 333: 	965 
    -- CP-element group 333:  members (22) 
      -- CP-element group 333: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588__exit__
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682
      -- CP-element group 333: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/$exit
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2591/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2601/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2601/SplitProtocol/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2601/SplitProtocol/Sample/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2601/SplitProtocol/Sample/rr
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2601/SplitProtocol/Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2601/SplitProtocol/Update/cr
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Sample/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Sample/rr
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Update/cr
      -- 
    rr_12315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(333), ack => type_cast_2601_inst_req_0); -- 
    cr_12320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(333), ack => type_cast_2601_inst_req_1); -- 
    rr_12338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(333), ack => type_cast_2607_inst_req_0); -- 
    cr_12343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(333), ack => type_cast_2607_inst_req_1); -- 
    zeropad3D_cp_element_group_333: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_333"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(318) & zeropad3D_CP_2152_elements(320) & zeropad3D_CP_2152_elements(326) & zeropad3D_CP_2152_elements(328) & zeropad3D_CP_2152_elements(330) & zeropad3D_CP_2152_elements(332);
      gj_zeropad3D_cp_element_group_333 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(333), clk => clk, reset => reset); --
    end block;
    -- CP-element group 334:  transition  input  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	972 
    -- CP-element group 334: successors 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/type_cast_2614_sample_completed_
      -- CP-element group 334: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/type_cast_2614_Sample/$exit
      -- CP-element group 334: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/type_cast_2614_Sample/ra
      -- 
    ra_6169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2614_inst_ack_0, ack => zeropad3D_CP_2152_elements(334)); -- 
    -- CP-element group 335:  branch  transition  place  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	972 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335: 	337 
    -- CP-element group 335:  members (13) 
      -- CP-element group 335: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622__exit__
      -- CP-element group 335: 	 branch_block_stmt_714/if_stmt_2623__entry__
      -- CP-element group 335: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/$exit
      -- CP-element group 335: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/type_cast_2614_update_completed_
      -- CP-element group 335: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/type_cast_2614_Update/$exit
      -- CP-element group 335: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/type_cast_2614_Update/ca
      -- CP-element group 335: 	 branch_block_stmt_714/if_stmt_2623_dead_link/$entry
      -- CP-element group 335: 	 branch_block_stmt_714/if_stmt_2623_eval_test/$entry
      -- CP-element group 335: 	 branch_block_stmt_714/if_stmt_2623_eval_test/$exit
      -- CP-element group 335: 	 branch_block_stmt_714/if_stmt_2623_eval_test/branch_req
      -- CP-element group 335: 	 branch_block_stmt_714/R_cmp687_2624_place
      -- CP-element group 335: 	 branch_block_stmt_714/if_stmt_2623_if_link/$entry
      -- CP-element group 335: 	 branch_block_stmt_714/if_stmt_2623_else_link/$entry
      -- 
    ca_6174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2614_inst_ack_1, ack => zeropad3D_CP_2152_elements(335)); -- 
    branch_req_6182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(335), ack => if_stmt_2623_branch_req_0); -- 
    -- CP-element group 336:  transition  place  input  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	973 
    -- CP-element group 336:  members (5) 
      -- CP-element group 336: 	 branch_block_stmt_714/if_stmt_2623_if_link/$exit
      -- CP-element group 336: 	 branch_block_stmt_714/if_stmt_2623_if_link/if_choice_transition
      -- CP-element group 336: 	 branch_block_stmt_714/whilex_xbody682_ifx_xthen717
      -- CP-element group 336: 	 branch_block_stmt_714/whilex_xbody682_ifx_xthen717_PhiReq/$entry
      -- CP-element group 336: 	 branch_block_stmt_714/whilex_xbody682_ifx_xthen717_PhiReq/$exit
      -- 
    if_choice_transition_6187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2623_branch_ack_1, ack => zeropad3D_CP_2152_elements(336)); -- 
    -- CP-element group 337:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337: 	339 
    -- CP-element group 337: 	341 
    -- CP-element group 337:  members (27) 
      -- CP-element group 337: 	 branch_block_stmt_714/merge_stmt_2629__exit__
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654__entry__
      -- CP-element group 337: 	 branch_block_stmt_714/if_stmt_2623_else_link/$exit
      -- CP-element group 337: 	 branch_block_stmt_714/if_stmt_2623_else_link/else_choice_transition
      -- CP-element group 337: 	 branch_block_stmt_714/whilex_xbody682_lorx_xlhsx_xfalse689
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/$entry
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_update_start_
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_word_address_calculated
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_root_address_calculated
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Sample/word_access_start/$entry
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Sample/word_access_start/word_0/$entry
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Sample/word_access_start/word_0/rr
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Update/word_access_complete/$entry
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Update/word_access_complete/word_0/$entry
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Update/word_access_complete/word_0/cr
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/type_cast_2635_update_start_
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/type_cast_2635_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/type_cast_2635_Update/cr
      -- CP-element group 337: 	 branch_block_stmt_714/whilex_xbody682_lorx_xlhsx_xfalse689_PhiReq/$entry
      -- CP-element group 337: 	 branch_block_stmt_714/whilex_xbody682_lorx_xlhsx_xfalse689_PhiReq/$exit
      -- CP-element group 337: 	 branch_block_stmt_714/merge_stmt_2629_PhiReqMerge
      -- CP-element group 337: 	 branch_block_stmt_714/merge_stmt_2629_PhiAck/$entry
      -- CP-element group 337: 	 branch_block_stmt_714/merge_stmt_2629_PhiAck/$exit
      -- CP-element group 337: 	 branch_block_stmt_714/merge_stmt_2629_PhiAck/dummy
      -- 
    else_choice_transition_6191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2623_branch_ack_0, ack => zeropad3D_CP_2152_elements(337)); -- 
    rr_6212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(337), ack => LOAD_row_high_2631_load_0_req_0); -- 
    cr_6223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(337), ack => LOAD_row_high_2631_load_0_req_1); -- 
    cr_6242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(337), ack => type_cast_2635_inst_req_1); -- 
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338:  members (5) 
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_sample_completed_
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Sample/$exit
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Sample/word_access_start/$exit
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Sample/word_access_start/word_0/$exit
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Sample/word_access_start/word_0/ra
      -- 
    ra_6213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2631_load_0_ack_0, ack => zeropad3D_CP_2152_elements(338)); -- 
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	337 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (12) 
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_update_completed_
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Update/$exit
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Update/word_access_complete/$exit
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Update/word_access_complete/word_0/$exit
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Update/word_access_complete/word_0/ca
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Update/LOAD_row_high_2631_Merge/$entry
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Update/LOAD_row_high_2631_Merge/$exit
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Update/LOAD_row_high_2631_Merge/merge_req
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/LOAD_row_high_2631_Update/LOAD_row_high_2631_Merge/merge_ack
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/type_cast_2635_sample_start_
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/type_cast_2635_Sample/$entry
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/type_cast_2635_Sample/rr
      -- 
    ca_6224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2631_load_0_ack_1, ack => zeropad3D_CP_2152_elements(339)); -- 
    rr_6237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(339), ack => type_cast_2635_inst_req_0); -- 
    -- CP-element group 340:  transition  input  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/type_cast_2635_sample_completed_
      -- CP-element group 340: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/type_cast_2635_Sample/$exit
      -- CP-element group 340: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/type_cast_2635_Sample/ra
      -- 
    ra_6238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2635_inst_ack_0, ack => zeropad3D_CP_2152_elements(340)); -- 
    -- CP-element group 341:  branch  transition  place  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	337 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341: 	343 
    -- CP-element group 341:  members (13) 
      -- CP-element group 341: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654__exit__
      -- CP-element group 341: 	 branch_block_stmt_714/if_stmt_2655__entry__
      -- CP-element group 341: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/$exit
      -- CP-element group 341: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/type_cast_2635_update_completed_
      -- CP-element group 341: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/type_cast_2635_Update/$exit
      -- CP-element group 341: 	 branch_block_stmt_714/assign_stmt_2632_to_assign_stmt_2654/type_cast_2635_Update/ca
      -- CP-element group 341: 	 branch_block_stmt_714/if_stmt_2655_dead_link/$entry
      -- CP-element group 341: 	 branch_block_stmt_714/if_stmt_2655_eval_test/$entry
      -- CP-element group 341: 	 branch_block_stmt_714/if_stmt_2655_eval_test/$exit
      -- CP-element group 341: 	 branch_block_stmt_714/if_stmt_2655_eval_test/branch_req
      -- CP-element group 341: 	 branch_block_stmt_714/R_cmp698_2656_place
      -- CP-element group 341: 	 branch_block_stmt_714/if_stmt_2655_if_link/$entry
      -- CP-element group 341: 	 branch_block_stmt_714/if_stmt_2655_else_link/$entry
      -- 
    ca_6243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2635_inst_ack_1, ack => zeropad3D_CP_2152_elements(341)); -- 
    branch_req_6251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(341), ack => if_stmt_2655_branch_req_0); -- 
    -- CP-element group 342:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342: 	345 
    -- CP-element group 342:  members (18) 
      -- CP-element group 342: 	 branch_block_stmt_714/merge_stmt_2661__exit__
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673__entry__
      -- CP-element group 342: 	 branch_block_stmt_714/if_stmt_2655_if_link/$exit
      -- CP-element group 342: 	 branch_block_stmt_714/if_stmt_2655_if_link/if_choice_transition
      -- CP-element group 342: 	 branch_block_stmt_714/lorx_xlhsx_xfalse689_lorx_xlhsx_xfalse700
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/$entry
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/type_cast_2665_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/type_cast_2665_update_start_
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/type_cast_2665_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/type_cast_2665_Sample/rr
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/type_cast_2665_Update/$entry
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/type_cast_2665_Update/cr
      -- CP-element group 342: 	 branch_block_stmt_714/lorx_xlhsx_xfalse689_lorx_xlhsx_xfalse700_PhiReq/$entry
      -- CP-element group 342: 	 branch_block_stmt_714/lorx_xlhsx_xfalse689_lorx_xlhsx_xfalse700_PhiReq/$exit
      -- CP-element group 342: 	 branch_block_stmt_714/merge_stmt_2661_PhiReqMerge
      -- CP-element group 342: 	 branch_block_stmt_714/merge_stmt_2661_PhiAck/$entry
      -- CP-element group 342: 	 branch_block_stmt_714/merge_stmt_2661_PhiAck/$exit
      -- CP-element group 342: 	 branch_block_stmt_714/merge_stmt_2661_PhiAck/dummy
      -- 
    if_choice_transition_6256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2655_branch_ack_1, ack => zeropad3D_CP_2152_elements(342)); -- 
    rr_6273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(342), ack => type_cast_2665_inst_req_0); -- 
    cr_6278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(342), ack => type_cast_2665_inst_req_1); -- 
    -- CP-element group 343:  transition  place  input  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	341 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	973 
    -- CP-element group 343:  members (5) 
      -- CP-element group 343: 	 branch_block_stmt_714/if_stmt_2655_else_link/$exit
      -- CP-element group 343: 	 branch_block_stmt_714/if_stmt_2655_else_link/else_choice_transition
      -- CP-element group 343: 	 branch_block_stmt_714/lorx_xlhsx_xfalse689_ifx_xthen717
      -- CP-element group 343: 	 branch_block_stmt_714/lorx_xlhsx_xfalse689_ifx_xthen717_PhiReq/$entry
      -- CP-element group 343: 	 branch_block_stmt_714/lorx_xlhsx_xfalse689_ifx_xthen717_PhiReq/$exit
      -- 
    else_choice_transition_6260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2655_branch_ack_0, ack => zeropad3D_CP_2152_elements(343)); -- 
    -- CP-element group 344:  transition  input  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: successors 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/type_cast_2665_sample_completed_
      -- CP-element group 344: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/type_cast_2665_Sample/$exit
      -- CP-element group 344: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/type_cast_2665_Sample/ra
      -- 
    ra_6274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2665_inst_ack_0, ack => zeropad3D_CP_2152_elements(344)); -- 
    -- CP-element group 345:  branch  transition  place  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	342 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (13) 
      -- CP-element group 345: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673__exit__
      -- CP-element group 345: 	 branch_block_stmt_714/if_stmt_2674__entry__
      -- CP-element group 345: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/$exit
      -- CP-element group 345: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/type_cast_2665_update_completed_
      -- CP-element group 345: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/type_cast_2665_Update/$exit
      -- CP-element group 345: 	 branch_block_stmt_714/assign_stmt_2666_to_assign_stmt_2673/type_cast_2665_Update/ca
      -- CP-element group 345: 	 branch_block_stmt_714/if_stmt_2674_dead_link/$entry
      -- CP-element group 345: 	 branch_block_stmt_714/if_stmt_2674_eval_test/$entry
      -- CP-element group 345: 	 branch_block_stmt_714/if_stmt_2674_eval_test/$exit
      -- CP-element group 345: 	 branch_block_stmt_714/if_stmt_2674_eval_test/branch_req
      -- CP-element group 345: 	 branch_block_stmt_714/R_cmp705_2675_place
      -- CP-element group 345: 	 branch_block_stmt_714/if_stmt_2674_if_link/$entry
      -- CP-element group 345: 	 branch_block_stmt_714/if_stmt_2674_else_link/$entry
      -- 
    ca_6279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2665_inst_ack_1, ack => zeropad3D_CP_2152_elements(345)); -- 
    branch_req_6287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(345), ack => if_stmt_2674_branch_req_0); -- 
    -- CP-element group 346:  transition  place  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	973 
    -- CP-element group 346:  members (5) 
      -- CP-element group 346: 	 branch_block_stmt_714/if_stmt_2674_if_link/$exit
      -- CP-element group 346: 	 branch_block_stmt_714/if_stmt_2674_if_link/if_choice_transition
      -- CP-element group 346: 	 branch_block_stmt_714/lorx_xlhsx_xfalse700_ifx_xthen717
      -- CP-element group 346: 	 branch_block_stmt_714/lorx_xlhsx_xfalse700_ifx_xthen717_PhiReq/$entry
      -- CP-element group 346: 	 branch_block_stmt_714/lorx_xlhsx_xfalse700_ifx_xthen717_PhiReq/$exit
      -- 
    if_choice_transition_6292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2674_branch_ack_1, ack => zeropad3D_CP_2152_elements(346)); -- 
    -- CP-element group 347:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347: 	349 
    -- CP-element group 347: 	351 
    -- CP-element group 347:  members (27) 
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699__entry__
      -- CP-element group 347: 	 branch_block_stmt_714/merge_stmt_2680__exit__
      -- CP-element group 347: 	 branch_block_stmt_714/if_stmt_2674_else_link/$exit
      -- CP-element group 347: 	 branch_block_stmt_714/if_stmt_2674_else_link/else_choice_transition
      -- CP-element group 347: 	 branch_block_stmt_714/lorx_xlhsx_xfalse700_lorx_xlhsx_xfalse707
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/$entry
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_sample_start_
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_update_start_
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_word_address_calculated
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_root_address_calculated
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Sample/$entry
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Sample/word_access_start/$entry
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Sample/word_access_start/word_0/$entry
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Sample/word_access_start/word_0/rr
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Update/word_access_complete/$entry
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Update/word_access_complete/word_0/$entry
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Update/word_access_complete/word_0/cr
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/type_cast_2686_update_start_
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/type_cast_2686_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/type_cast_2686_Update/cr
      -- CP-element group 347: 	 branch_block_stmt_714/lorx_xlhsx_xfalse700_lorx_xlhsx_xfalse707_PhiReq/$entry
      -- CP-element group 347: 	 branch_block_stmt_714/lorx_xlhsx_xfalse700_lorx_xlhsx_xfalse707_PhiReq/$exit
      -- CP-element group 347: 	 branch_block_stmt_714/merge_stmt_2680_PhiReqMerge
      -- CP-element group 347: 	 branch_block_stmt_714/merge_stmt_2680_PhiAck/$entry
      -- CP-element group 347: 	 branch_block_stmt_714/merge_stmt_2680_PhiAck/$exit
      -- CP-element group 347: 	 branch_block_stmt_714/merge_stmt_2680_PhiAck/dummy
      -- 
    else_choice_transition_6296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2674_branch_ack_0, ack => zeropad3D_CP_2152_elements(347)); -- 
    rr_6317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(347), ack => LOAD_col_high_2682_load_0_req_0); -- 
    cr_6328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(347), ack => LOAD_col_high_2682_load_0_req_1); -- 
    cr_6347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(347), ack => type_cast_2686_inst_req_1); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348:  members (5) 
      -- CP-element group 348: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_sample_completed_
      -- CP-element group 348: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Sample/$exit
      -- CP-element group 348: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Sample/word_access_start/$exit
      -- CP-element group 348: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Sample/word_access_start/word_0/$exit
      -- CP-element group 348: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Sample/word_access_start/word_0/ra
      -- 
    ra_6318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2682_load_0_ack_0, ack => zeropad3D_CP_2152_elements(348)); -- 
    -- CP-element group 349:  transition  input  output  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	347 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	350 
    -- CP-element group 349:  members (12) 
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_update_completed_
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Update/$exit
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Update/word_access_complete/$exit
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Update/word_access_complete/word_0/$exit
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Update/word_access_complete/word_0/ca
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Update/LOAD_col_high_2682_Merge/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Update/LOAD_col_high_2682_Merge/$exit
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Update/LOAD_col_high_2682_Merge/merge_req
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/LOAD_col_high_2682_Update/LOAD_col_high_2682_Merge/merge_ack
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/type_cast_2686_sample_start_
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/type_cast_2686_Sample/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/type_cast_2686_Sample/rr
      -- 
    ca_6329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2682_load_0_ack_1, ack => zeropad3D_CP_2152_elements(349)); -- 
    rr_6342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(349), ack => type_cast_2686_inst_req_0); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	349 
    -- CP-element group 350: successors 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/type_cast_2686_sample_completed_
      -- CP-element group 350: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/type_cast_2686_Sample/$exit
      -- CP-element group 350: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/type_cast_2686_Sample/ra
      -- 
    ra_6343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2686_inst_ack_0, ack => zeropad3D_CP_2152_elements(350)); -- 
    -- CP-element group 351:  branch  transition  place  input  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	347 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351: 	353 
    -- CP-element group 351:  members (13) 
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2700__entry__
      -- CP-element group 351: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699__exit__
      -- CP-element group 351: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/$exit
      -- CP-element group 351: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/type_cast_2686_update_completed_
      -- CP-element group 351: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/type_cast_2686_Update/$exit
      -- CP-element group 351: 	 branch_block_stmt_714/assign_stmt_2683_to_assign_stmt_2699/type_cast_2686_Update/ca
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2700_dead_link/$entry
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2700_eval_test/$entry
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2700_eval_test/$exit
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2700_eval_test/branch_req
      -- CP-element group 351: 	 branch_block_stmt_714/R_cmp715_2701_place
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2700_if_link/$entry
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2700_else_link/$entry
      -- 
    ca_6348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2686_inst_ack_1, ack => zeropad3D_CP_2152_elements(351)); -- 
    branch_req_6356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(351), ack => if_stmt_2700_branch_req_0); -- 
    -- CP-element group 352:  fork  transition  place  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	368 
    -- CP-element group 352: 	369 
    -- CP-element group 352: 	371 
    -- CP-element group 352: 	373 
    -- CP-element group 352: 	375 
    -- CP-element group 352: 	377 
    -- CP-element group 352: 	379 
    -- CP-element group 352: 	381 
    -- CP-element group 352: 	383 
    -- CP-element group 352: 	386 
    -- CP-element group 352:  members (46) 
      -- CP-element group 352: 	 branch_block_stmt_714/merge_stmt_2764__exit__
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869__entry__
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2857_update_start_
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2857_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_final_index_sum_regn_update_start
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Update/word_access_complete/word_0/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_update_start_
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Update/word_access_complete/word_0/cr
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Update/word_access_complete/word_0/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Update/word_access_complete/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2864_complete/req
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_final_index_sum_regn_Update/req
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Update/word_access_complete/word_0/cr
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_final_index_sum_regn_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2864_update_start_
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2857_Update/cr
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2864_complete/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Update/word_access_complete/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/if_stmt_2700_if_link/$exit
      -- CP-element group 352: 	 branch_block_stmt_714/if_stmt_2700_if_link/if_choice_transition
      -- CP-element group 352: 	 branch_block_stmt_714/lorx_xlhsx_xfalse707_ifx_xelse738
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2768_sample_start_
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2768_update_start_
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2768_Sample/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2768_Sample/rr
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2768_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2768_Update/cr
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2832_update_start_
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2832_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2832_Update/cr
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2839_update_start_
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_final_index_sum_regn_update_start
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_final_index_sum_regn_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_final_index_sum_regn_Update/req
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2839_complete/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2839_complete/req
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_update_start_
      -- CP-element group 352: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/lorx_xlhsx_xfalse707_ifx_xelse738_PhiReq/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/lorx_xlhsx_xfalse707_ifx_xelse738_PhiReq/$exit
      -- CP-element group 352: 	 branch_block_stmt_714/merge_stmt_2764_PhiReqMerge
      -- CP-element group 352: 	 branch_block_stmt_714/merge_stmt_2764_PhiAck/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/merge_stmt_2764_PhiAck/$exit
      -- CP-element group 352: 	 branch_block_stmt_714/merge_stmt_2764_PhiAck/dummy
      -- 
    if_choice_transition_6361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2700_branch_ack_1, ack => zeropad3D_CP_2152_elements(352)); -- 
    cr_6744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(352), ack => ptr_deref_2867_store_0_req_1); -- 
    req_6694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(352), ack => addr_of_2864_final_reg_req_1); -- 
    req_6679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(352), ack => array_obj_ref_2863_index_offset_req_1); -- 
    cr_6629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(352), ack => ptr_deref_2843_load_0_req_1); -- 
    cr_6648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(352), ack => type_cast_2857_inst_req_1); -- 
    rr_6519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(352), ack => type_cast_2768_inst_req_0); -- 
    cr_6524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(352), ack => type_cast_2768_inst_req_1); -- 
    cr_6538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(352), ack => type_cast_2832_inst_req_1); -- 
    req_6569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(352), ack => array_obj_ref_2838_index_offset_req_1); -- 
    req_6584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(352), ack => addr_of_2839_final_reg_req_1); -- 
    -- CP-element group 353:  transition  place  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	351 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	973 
    -- CP-element group 353:  members (5) 
      -- CP-element group 353: 	 branch_block_stmt_714/if_stmt_2700_else_link/$exit
      -- CP-element group 353: 	 branch_block_stmt_714/if_stmt_2700_else_link/else_choice_transition
      -- CP-element group 353: 	 branch_block_stmt_714/lorx_xlhsx_xfalse707_ifx_xthen717
      -- CP-element group 353: 	 branch_block_stmt_714/lorx_xlhsx_xfalse707_ifx_xthen717_PhiReq/$entry
      -- CP-element group 353: 	 branch_block_stmt_714/lorx_xlhsx_xfalse707_ifx_xthen717_PhiReq/$exit
      -- 
    else_choice_transition_6365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2700_branch_ack_0, ack => zeropad3D_CP_2152_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	973 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2710_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2710_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2710_Sample/ra
      -- 
    ra_6379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2710_inst_ack_0, ack => zeropad3D_CP_2152_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	973 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	358 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2710_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2710_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2710_Update/ca
      -- 
    ca_6384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2710_inst_ack_1, ack => zeropad3D_CP_2152_elements(355)); -- 
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	973 
    -- CP-element group 356: successors 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2715_sample_completed_
      -- CP-element group 356: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2715_Sample/$exit
      -- CP-element group 356: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2715_Sample/ra
      -- 
    ra_6393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2715_inst_ack_0, ack => zeropad3D_CP_2152_elements(356)); -- 
    -- CP-element group 357:  transition  input  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	973 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2715_update_completed_
      -- CP-element group 357: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2715_Update/$exit
      -- CP-element group 357: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2715_Update/ca
      -- 
    ca_6398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2715_inst_ack_1, ack => zeropad3D_CP_2152_elements(357)); -- 
    -- CP-element group 358:  join  transition  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	355 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2749_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2749_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2749_Sample/rr
      -- 
    rr_6406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(358), ack => type_cast_2749_inst_req_0); -- 
    zeropad3D_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(355) & zeropad3D_CP_2152_elements(357);
      gj_zeropad3D_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  transition  input  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2749_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2749_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2749_Sample/ra
      -- 
    ra_6407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2749_inst_ack_0, ack => zeropad3D_CP_2152_elements(359)); -- 
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	973 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (16) 
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2749_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2749_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2749_Update/ca
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_index_resized_1
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_index_scaled_1
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_index_computed_1
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_index_resize_1/$entry
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_index_resize_1/$exit
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_index_resize_1/index_resize_req
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_index_resize_1/index_resize_ack
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_index_scale_1/$entry
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_index_scale_1/$exit
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_index_scale_1/scale_rename_req
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_index_scale_1/scale_rename_ack
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_final_index_sum_regn_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_final_index_sum_regn_Sample/req
      -- 
    ca_6412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2749_inst_ack_1, ack => zeropad3D_CP_2152_elements(360)); -- 
    req_6437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(360), ack => array_obj_ref_2755_index_offset_req_0); -- 
    -- CP-element group 361:  transition  input  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	367 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_final_index_sum_regn_sample_complete
      -- CP-element group 361: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_final_index_sum_regn_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_final_index_sum_regn_Sample/ack
      -- 
    ack_6438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2755_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(361)); -- 
    -- CP-element group 362:  transition  input  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	973 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (11) 
      -- CP-element group 362: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/addr_of_2756_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_root_address_calculated
      -- CP-element group 362: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_offset_calculated
      -- CP-element group 362: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_final_index_sum_regn_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_final_index_sum_regn_Update/ack
      -- CP-element group 362: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_base_plus_offset/$entry
      -- CP-element group 362: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_base_plus_offset/$exit
      -- CP-element group 362: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_base_plus_offset/sum_rename_req
      -- CP-element group 362: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_base_plus_offset/sum_rename_ack
      -- CP-element group 362: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/addr_of_2756_request/$entry
      -- CP-element group 362: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/addr_of_2756_request/req
      -- 
    ack_6443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2755_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(362)); -- 
    req_6452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(362), ack => addr_of_2756_final_reg_req_0); -- 
    -- CP-element group 363:  transition  input  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/addr_of_2756_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/addr_of_2756_request/$exit
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/addr_of_2756_request/ack
      -- 
    ack_6453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2756_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(363)); -- 
    -- CP-element group 364:  join  fork  transition  input  output  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	973 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (28) 
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/addr_of_2756_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/addr_of_2756_complete/$exit
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/addr_of_2756_complete/ack
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_sample_start_
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_base_address_calculated
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_word_address_calculated
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_root_address_calculated
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_base_address_resized
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_base_addr_resize/$entry
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_base_addr_resize/$exit
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_base_addr_resize/base_resize_req
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_base_addr_resize/base_resize_ack
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_base_plus_offset/$entry
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_base_plus_offset/$exit
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_base_plus_offset/sum_rename_req
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_base_plus_offset/sum_rename_ack
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_word_addrgen/$entry
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_word_addrgen/$exit
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_word_addrgen/root_register_req
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_word_addrgen/root_register_ack
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Sample/$entry
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Sample/ptr_deref_2759_Split/$entry
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Sample/ptr_deref_2759_Split/$exit
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Sample/ptr_deref_2759_Split/split_req
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Sample/ptr_deref_2759_Split/split_ack
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Sample/word_access_start/$entry
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Sample/word_access_start/word_0/$entry
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Sample/word_access_start/word_0/rr
      -- 
    ack_6458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2756_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(364)); -- 
    rr_6496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(364), ack => ptr_deref_2759_store_0_req_0); -- 
    -- CP-element group 365:  transition  input  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365:  members (5) 
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Sample/word_access_start/$exit
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Sample/word_access_start/word_0/$exit
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Sample/word_access_start/word_0/ra
      -- 
    ra_6497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2759_store_0_ack_0, ack => zeropad3D_CP_2152_elements(365)); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	973 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366:  members (5) 
      -- CP-element group 366: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Update/word_access_complete/$exit
      -- CP-element group 366: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Update/word_access_complete/word_0/$exit
      -- CP-element group 366: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Update/word_access_complete/word_0/ca
      -- 
    ca_6508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2759_store_0_ack_1, ack => zeropad3D_CP_2152_elements(366)); -- 
    -- CP-element group 367:  join  transition  place  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	361 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	974 
    -- CP-element group 367:  members (5) 
      -- CP-element group 367: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762__exit__
      -- CP-element group 367: 	 branch_block_stmt_714/ifx_xthen717_ifx_xend786
      -- CP-element group 367: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/$exit
      -- CP-element group 367: 	 branch_block_stmt_714/ifx_xthen717_ifx_xend786_PhiReq/$entry
      -- CP-element group 367: 	 branch_block_stmt_714/ifx_xthen717_ifx_xend786_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_367: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_367"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(361) & zeropad3D_CP_2152_elements(366);
      gj_zeropad3D_cp_element_group_367 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	352 
    -- CP-element group 368: successors 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2768_sample_completed_
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2768_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2768_Sample/ra
      -- 
    ra_6520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2768_inst_ack_0, ack => zeropad3D_CP_2152_elements(368)); -- 
    -- CP-element group 369:  fork  transition  input  output  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	352 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369: 	378 
    -- CP-element group 369:  members (9) 
      -- CP-element group 369: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2857_sample_start_
      -- CP-element group 369: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2857_Sample/$entry
      -- CP-element group 369: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2857_Sample/rr
      -- CP-element group 369: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2768_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2768_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2768_Update/ca
      -- CP-element group 369: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2832_sample_start_
      -- CP-element group 369: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2832_Sample/$entry
      -- CP-element group 369: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2832_Sample/rr
      -- 
    ca_6525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2768_inst_ack_1, ack => zeropad3D_CP_2152_elements(369)); -- 
    rr_6533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(369), ack => type_cast_2832_inst_req_0); -- 
    rr_6643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(369), ack => type_cast_2857_inst_req_0); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2832_sample_completed_
      -- CP-element group 370: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2832_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2832_Sample/ra
      -- 
    ra_6534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2832_inst_ack_0, ack => zeropad3D_CP_2152_elements(370)); -- 
    -- CP-element group 371:  transition  input  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	352 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (16) 
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2832_update_completed_
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2832_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2832_Update/ca
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_index_resized_1
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_index_scaled_1
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_index_computed_1
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_index_resize_1/$entry
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_index_resize_1/$exit
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_index_resize_1/index_resize_req
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_index_resize_1/index_resize_ack
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_index_scale_1/$entry
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_index_scale_1/$exit
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_index_scale_1/scale_rename_req
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_index_scale_1/scale_rename_ack
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_final_index_sum_regn_Sample/$entry
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_final_index_sum_regn_Sample/req
      -- 
    ca_6539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2832_inst_ack_1, ack => zeropad3D_CP_2152_elements(371)); -- 
    req_6564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(371), ack => array_obj_ref_2838_index_offset_req_0); -- 
    -- CP-element group 372:  transition  input  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	387 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_final_index_sum_regn_sample_complete
      -- CP-element group 372: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_final_index_sum_regn_Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_final_index_sum_regn_Sample/ack
      -- 
    ack_6565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2838_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(372)); -- 
    -- CP-element group 373:  transition  input  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	352 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (11) 
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2839_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_root_address_calculated
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_offset_calculated
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_final_index_sum_regn_Update/$exit
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_final_index_sum_regn_Update/ack
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_base_plus_offset/$entry
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_base_plus_offset/$exit
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_base_plus_offset/sum_rename_req
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2838_base_plus_offset/sum_rename_ack
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2839_request/$entry
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2839_request/req
      -- 
    ack_6570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2838_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(373)); -- 
    req_6579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(373), ack => addr_of_2839_final_reg_req_0); -- 
    -- CP-element group 374:  transition  input  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2839_sample_completed_
      -- CP-element group 374: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2839_request/$exit
      -- CP-element group 374: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2839_request/ack
      -- 
    ack_6580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2839_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(374)); -- 
    -- CP-element group 375:  join  fork  transition  input  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	352 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (24) 
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2839_update_completed_
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2839_complete/$exit
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2839_complete/ack
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_base_address_calculated
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_word_address_calculated
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_root_address_calculated
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_base_address_resized
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_base_addr_resize/$entry
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_base_addr_resize/$exit
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_base_addr_resize/base_resize_req
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_base_addr_resize/base_resize_ack
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_base_plus_offset/$entry
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_base_plus_offset/$exit
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_base_plus_offset/sum_rename_req
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_base_plus_offset/sum_rename_ack
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_word_addrgen/$entry
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_word_addrgen/$exit
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_word_addrgen/root_register_req
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_word_addrgen/root_register_ack
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Sample/word_access_start/$entry
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Sample/word_access_start/word_0/$entry
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Sample/word_access_start/word_0/rr
      -- 
    ack_6585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2839_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(375)); -- 
    rr_6618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(375), ack => ptr_deref_2843_load_0_req_0); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376:  members (5) 
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_sample_completed_
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Sample/word_access_start/$exit
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Sample/word_access_start/word_0/$exit
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Sample/word_access_start/word_0/ra
      -- 
    ra_6619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2843_load_0_ack_0, ack => zeropad3D_CP_2152_elements(376)); -- 
    -- CP-element group 377:  transition  input  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	352 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	384 
    -- CP-element group 377:  members (9) 
      -- CP-element group 377: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Update/ptr_deref_2843_Merge/merge_ack
      -- CP-element group 377: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Update/ptr_deref_2843_Merge/merge_req
      -- CP-element group 377: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Update/ptr_deref_2843_Merge/$exit
      -- CP-element group 377: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Update/ptr_deref_2843_Merge/$entry
      -- CP-element group 377: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Update/word_access_complete/word_0/ca
      -- CP-element group 377: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Update/word_access_complete/word_0/$exit
      -- CP-element group 377: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Update/word_access_complete/$exit
      -- CP-element group 377: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_update_completed_
      -- CP-element group 377: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2843_Update/$exit
      -- 
    ca_6630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2843_load_0_ack_1, ack => zeropad3D_CP_2152_elements(377)); -- 
    -- CP-element group 378:  transition  input  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	369 
    -- CP-element group 378: successors 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2857_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2857_Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2857_Sample/ra
      -- 
    ra_6644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2857_inst_ack_0, ack => zeropad3D_CP_2152_elements(378)); -- 
    -- CP-element group 379:  transition  input  output  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	352 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379:  members (16) 
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_index_resize_1/$entry
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_index_resize_1/$exit
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_index_resize_1/index_resize_req
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_index_resize_1/index_resize_ack
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_index_scale_1/$entry
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2857_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_index_scale_1/$exit
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_index_scale_1/scale_rename_req
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_index_scale_1/scale_rename_ack
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_index_computed_1
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_index_scaled_1
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_index_resized_1
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2857_Update/ca
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_final_index_sum_regn_Sample/req
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_final_index_sum_regn_Sample/$entry
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/type_cast_2857_Update/$exit
      -- 
    ca_6649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2857_inst_ack_1, ack => zeropad3D_CP_2152_elements(379)); -- 
    req_6674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(379), ack => array_obj_ref_2863_index_offset_req_0); -- 
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	379 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	387 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_final_index_sum_regn_sample_complete
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_final_index_sum_regn_Sample/ack
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_final_index_sum_regn_Sample/$exit
      -- 
    ack_6675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2863_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(380)); -- 
    -- CP-element group 381:  transition  input  output  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	352 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (11) 
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2864_request/req
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2864_request/$entry
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_offset_calculated
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_root_address_calculated
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_base_plus_offset/sum_rename_ack
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_base_plus_offset/sum_rename_req
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_base_plus_offset/$exit
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_base_plus_offset/$entry
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_final_index_sum_regn_Update/ack
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/array_obj_ref_2863_final_index_sum_regn_Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2864_sample_start_
      -- 
    ack_6680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2863_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(381)); -- 
    req_6689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(381), ack => addr_of_2864_final_reg_req_0); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2864_request/$exit
      -- CP-element group 382: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2864_request/ack
      -- CP-element group 382: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2864_sample_completed_
      -- 
    ack_6690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2864_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(382)); -- 
    -- CP-element group 383:  fork  transition  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	352 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (19) 
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_base_addr_resize/$entry
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_base_addr_resize/$exit
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_base_addr_resize/base_resize_req
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_base_addr_resize/base_resize_ack
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_base_address_resized
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_root_address_calculated
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_word_address_calculated
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_base_address_calculated
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2864_update_completed_
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2864_complete/ack
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/addr_of_2864_complete/$exit
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_word_addrgen/root_register_ack
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_word_addrgen/root_register_req
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_word_addrgen/$exit
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_word_addrgen/$entry
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_base_plus_offset/sum_rename_ack
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_base_plus_offset/sum_rename_req
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_base_plus_offset/$exit
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_base_plus_offset/$entry
      -- 
    ack_6695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2864_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(383)); -- 
    -- CP-element group 384:  join  transition  output  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	377 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384:  members (9) 
      -- CP-element group 384: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_sample_start_
      -- CP-element group 384: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Sample/word_access_start/word_0/rr
      -- CP-element group 384: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Sample/word_access_start/word_0/$entry
      -- CP-element group 384: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Sample/word_access_start/$entry
      -- CP-element group 384: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Sample/ptr_deref_2867_Split/split_ack
      -- CP-element group 384: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Sample/ptr_deref_2867_Split/split_req
      -- CP-element group 384: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Sample/ptr_deref_2867_Split/$exit
      -- CP-element group 384: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Sample/ptr_deref_2867_Split/$entry
      -- CP-element group 384: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Sample/$entry
      -- 
    rr_6733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(384), ack => ptr_deref_2867_store_0_req_0); -- 
    zeropad3D_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(377) & zeropad3D_CP_2152_elements(383);
      gj_zeropad3D_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385:  members (5) 
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_sample_completed_
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Sample/word_access_start/word_0/ra
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Sample/word_access_start/word_0/$exit
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Sample/word_access_start/$exit
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Sample/$exit
      -- 
    ra_6734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2867_store_0_ack_0, ack => zeropad3D_CP_2152_elements(385)); -- 
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	352 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	387 
    -- CP-element group 386:  members (5) 
      -- CP-element group 386: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_update_completed_
      -- CP-element group 386: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Update/word_access_complete/word_0/ca
      -- CP-element group 386: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Update/word_access_complete/word_0/$exit
      -- CP-element group 386: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Update/word_access_complete/$exit
      -- CP-element group 386: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/ptr_deref_2867_Update/$exit
      -- 
    ca_6745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2867_store_0_ack_1, ack => zeropad3D_CP_2152_elements(386)); -- 
    -- CP-element group 387:  join  transition  place  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	372 
    -- CP-element group 387: 	380 
    -- CP-element group 387: 	386 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	974 
    -- CP-element group 387:  members (5) 
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869__exit__
      -- CP-element group 387: 	 branch_block_stmt_714/ifx_xelse738_ifx_xend786
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2769_to_assign_stmt_2869/$exit
      -- CP-element group 387: 	 branch_block_stmt_714/ifx_xelse738_ifx_xend786_PhiReq/$entry
      -- CP-element group 387: 	 branch_block_stmt_714/ifx_xelse738_ifx_xend786_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_387: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_387"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(372) & zeropad3D_CP_2152_elements(380) & zeropad3D_CP_2152_elements(386);
      gj_zeropad3D_cp_element_group_387 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(387), clk => clk, reset => reset); --
    end block;
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	974 
    -- CP-element group 388: successors 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/type_cast_2875_Sample/ra
      -- CP-element group 388: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/type_cast_2875_Sample/$exit
      -- CP-element group 388: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/type_cast_2875_sample_completed_
      -- 
    ra_6757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2875_inst_ack_0, ack => zeropad3D_CP_2152_elements(388)); -- 
    -- CP-element group 389:  branch  transition  place  input  output  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	974 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	390 
    -- CP-element group 389: 	391 
    -- CP-element group 389:  members (13) 
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889__exit__
      -- CP-element group 389: 	 branch_block_stmt_714/if_stmt_2890__entry__
      -- CP-element group 389: 	 branch_block_stmt_714/if_stmt_2890_else_link/$entry
      -- CP-element group 389: 	 branch_block_stmt_714/if_stmt_2890_if_link/$entry
      -- CP-element group 389: 	 branch_block_stmt_714/if_stmt_2890_eval_test/branch_req
      -- CP-element group 389: 	 branch_block_stmt_714/if_stmt_2890_eval_test/$exit
      -- CP-element group 389: 	 branch_block_stmt_714/if_stmt_2890_eval_test/$entry
      -- CP-element group 389: 	 branch_block_stmt_714/if_stmt_2890_dead_link/$entry
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/type_cast_2875_Update/ca
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/type_cast_2875_Update/$exit
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/type_cast_2875_update_completed_
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/$exit
      -- CP-element group 389: 	 branch_block_stmt_714/R_cmp794_2891_place
      -- 
    ca_6762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2875_inst_ack_1, ack => zeropad3D_CP_2152_elements(389)); -- 
    branch_req_6770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(389), ack => if_stmt_2890_branch_req_0); -- 
    -- CP-element group 390:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	389 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	983 
    -- CP-element group 390: 	984 
    -- CP-element group 390: 	986 
    -- CP-element group 390: 	987 
    -- CP-element group 390: 	989 
    -- CP-element group 390: 	990 
    -- CP-element group 390:  members (40) 
      -- CP-element group 390: 	 branch_block_stmt_714/merge_stmt_2896__exit__
      -- CP-element group 390: 	 branch_block_stmt_714/assign_stmt_2902__entry__
      -- CP-element group 390: 	 branch_block_stmt_714/assign_stmt_2902__exit__
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837
      -- CP-element group 390: 	 branch_block_stmt_714/assign_stmt_2902/$exit
      -- CP-element group 390: 	 branch_block_stmt_714/assign_stmt_2902/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/if_stmt_2890_if_link/if_choice_transition
      -- CP-element group 390: 	 branch_block_stmt_714/if_stmt_2890_if_link/$exit
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xend786_ifx_xthen796
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/type_cast_2986/SplitProtocol/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/type_cast_2986/SplitProtocol/Sample/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/type_cast_2986/SplitProtocol/Sample/rr
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/type_cast_2986/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/merge_stmt_2896_PhiReqMerge
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/merge_stmt_2896_PhiAck/dummy
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_2999/SplitProtocol/Update/cr
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_2999/SplitProtocol/Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_2999/SplitProtocol/Sample/rr
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_2999/SplitProtocol/Sample/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_2999/SplitProtocol/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/type_cast_2986/SplitProtocol/Update/cr
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_2999/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/type_cast_2986/SplitProtocol/Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/cr
      -- CP-element group 390: 	 branch_block_stmt_714/merge_stmt_2896_PhiAck/$exit
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/merge_stmt_2896_PhiAck/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/rr
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xend786_ifx_xthen796_PhiReq/$entry
      -- CP-element group 390: 	 branch_block_stmt_714/ifx_xend786_ifx_xthen796_PhiReq/$exit
      -- 
    if_choice_transition_6775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2890_branch_ack_1, ack => zeropad3D_CP_2152_elements(390)); -- 
    rr_12528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(390), ack => type_cast_2986_inst_req_0); -- 
    cr_12579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(390), ack => type_cast_2999_inst_req_1); -- 
    rr_12574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(390), ack => type_cast_2999_inst_req_0); -- 
    cr_12533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(390), ack => type_cast_2986_inst_req_1); -- 
    cr_12556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(390), ack => type_cast_2993_inst_req_1); -- 
    rr_12551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(390), ack => type_cast_2993_inst_req_0); -- 
    -- CP-element group 391:  fork  transition  place  input  output  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	389 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391: 	393 
    -- CP-element group 391: 	394 
    -- CP-element group 391: 	395 
    -- CP-element group 391: 	397 
    -- CP-element group 391: 	400 
    -- CP-element group 391: 	402 
    -- CP-element group 391: 	403 
    -- CP-element group 391: 	404 
    -- CP-element group 391: 	406 
    -- CP-element group 391:  members (54) 
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975__entry__
      -- CP-element group 391: 	 branch_block_stmt_714/merge_stmt_2904__exit__
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2914_update_start_
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2951_update_start_
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Sample/word_access_start/word_0/rr
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_word_address_calculated
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_root_address_calculated
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2914_Sample/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2921_Update/cr
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Sample/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2914_Sample/rr
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2914_Update/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2914_Update/cr
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Sample/word_access_start/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2935_update_start_
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Sample/word_access_start/word_0/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2935_Update/cr
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2914_sample_start_
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Sample/word_access_start/word_0/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2921_Update/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Update/word_access_complete/word_0/cr
      -- CP-element group 391: 	 branch_block_stmt_714/if_stmt_2890_else_link/else_choice_transition
      -- CP-element group 391: 	 branch_block_stmt_714/if_stmt_2890_else_link/$exit
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Update/word_access_complete/word_0/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Update/word_access_complete/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Sample/word_access_start/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2935_Update/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2951_Update/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2921_update_start_
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Sample/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_root_address_calculated
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_word_address_calculated
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Update/word_access_complete/word_0/cr
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Update/word_access_complete/word_0/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/ifx_xend786_ifx_xelse801
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_update_start_
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Update/word_access_complete/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_update_start_
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_sample_start_
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Update/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Update/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_sample_start_
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Sample/word_access_start/word_0/rr
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2951_Update/cr
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2958_update_start_
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2958_Update/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2958_Update/cr
      -- CP-element group 391: 	 branch_block_stmt_714/merge_stmt_2904_PhiReqMerge
      -- CP-element group 391: 	 branch_block_stmt_714/merge_stmt_2904_PhiAck/dummy
      -- CP-element group 391: 	 branch_block_stmt_714/merge_stmt_2904_PhiAck/$exit
      -- CP-element group 391: 	 branch_block_stmt_714/merge_stmt_2904_PhiAck/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/ifx_xend786_ifx_xelse801_PhiReq/$exit
      -- CP-element group 391: 	 branch_block_stmt_714/ifx_xend786_ifx_xelse801_PhiReq/$entry
      -- 
    else_choice_transition_6779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2890_branch_ack_0, ack => zeropad3D_CP_2152_elements(391)); -- 
    rr_6892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(391), ack => LOAD_row_high_2954_load_0_req_0); -- 
    cr_6847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(391), ack => type_cast_2921_inst_req_1); -- 
    rr_6795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(391), ack => type_cast_2914_inst_req_0); -- 
    cr_6800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(391), ack => type_cast_2914_inst_req_1); -- 
    cr_6861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(391), ack => type_cast_2935_inst_req_1); -- 
    cr_6903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(391), ack => LOAD_row_high_2954_load_0_req_1); -- 
    cr_6828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(391), ack => LOAD_col_high_2917_load_0_req_1); -- 
    rr_6817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(391), ack => LOAD_col_high_2917_load_0_req_0); -- 
    cr_6875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(391), ack => type_cast_2951_inst_req_1); -- 
    cr_6922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(391), ack => type_cast_2958_inst_req_1); -- 
    -- CP-element group 392:  transition  input  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	391 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2914_sample_completed_
      -- CP-element group 392: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2914_Sample/$exit
      -- CP-element group 392: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2914_Sample/ra
      -- 
    ra_6796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2914_inst_ack_0, ack => zeropad3D_CP_2152_elements(392)); -- 
    -- CP-element group 393:  transition  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	391 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	398 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2914_update_completed_
      -- CP-element group 393: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2914_Update/$exit
      -- CP-element group 393: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2914_Update/ca
      -- 
    ca_6801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2914_inst_ack_1, ack => zeropad3D_CP_2152_elements(393)); -- 
    -- CP-element group 394:  transition  input  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	391 
    -- CP-element group 394: successors 
    -- CP-element group 394:  members (5) 
      -- CP-element group 394: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Sample/$exit
      -- CP-element group 394: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Sample/word_access_start/$exit
      -- CP-element group 394: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Sample/word_access_start/word_0/$exit
      -- CP-element group 394: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_sample_completed_
      -- CP-element group 394: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Sample/word_access_start/word_0/ra
      -- 
    ra_6818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2917_load_0_ack_0, ack => zeropad3D_CP_2152_elements(394)); -- 
    -- CP-element group 395:  transition  input  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	391 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395:  members (12) 
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2921_Sample/rr
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2921_Sample/$entry
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2921_sample_start_
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Update/LOAD_col_high_2917_Merge/merge_ack
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Update/LOAD_col_high_2917_Merge/merge_req
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Update/LOAD_col_high_2917_Merge/$exit
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Update/LOAD_col_high_2917_Merge/$entry
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Update/word_access_complete/word_0/ca
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Update/word_access_complete/word_0/$exit
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Update/word_access_complete/$exit
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_update_completed_
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_col_high_2917_Update/$exit
      -- 
    ca_6829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2917_load_0_ack_1, ack => zeropad3D_CP_2152_elements(395)); -- 
    rr_6842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(395), ack => type_cast_2921_inst_req_0); -- 
    -- CP-element group 396:  transition  input  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2921_Sample/ra
      -- CP-element group 396: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2921_Sample/$exit
      -- CP-element group 396: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2921_sample_completed_
      -- 
    ra_6843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2921_inst_ack_0, ack => zeropad3D_CP_2152_elements(396)); -- 
    -- CP-element group 397:  transition  input  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	391 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2921_Update/$exit
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2921_Update/ca
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2921_update_completed_
      -- 
    ca_6848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2921_inst_ack_1, ack => zeropad3D_CP_2152_elements(397)); -- 
    -- CP-element group 398:  join  transition  output  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	393 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2935_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2935_Sample/rr
      -- CP-element group 398: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2935_Sample/$entry
      -- 
    rr_6856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(398), ack => type_cast_2935_inst_req_0); -- 
    zeropad3D_cp_element_group_398: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_398"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(393) & zeropad3D_CP_2152_elements(397);
      gj_zeropad3D_cp_element_group_398 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(398), clk => clk, reset => reset); --
    end block;
    -- CP-element group 399:  transition  input  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2935_sample_completed_
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2935_Sample/ra
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2935_Sample/$exit
      -- 
    ra_6857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2935_inst_ack_0, ack => zeropad3D_CP_2152_elements(399)); -- 
    -- CP-element group 400:  transition  input  output  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	391 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (6) 
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2951_Sample/$entry
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2935_update_completed_
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2951_sample_start_
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2935_Update/ca
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2935_Update/$exit
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2951_Sample/rr
      -- 
    ca_6862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2935_inst_ack_1, ack => zeropad3D_CP_2152_elements(400)); -- 
    rr_6870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(400), ack => type_cast_2951_inst_req_0); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2951_sample_completed_
      -- CP-element group 401: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2951_Sample/ra
      -- CP-element group 401: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2951_Sample/$exit
      -- 
    ra_6871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2951_inst_ack_0, ack => zeropad3D_CP_2152_elements(401)); -- 
    -- CP-element group 402:  transition  input  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	391 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	407 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2951_Update/$exit
      -- CP-element group 402: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2951_update_completed_
      -- CP-element group 402: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2951_Update/ca
      -- 
    ca_6876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2951_inst_ack_1, ack => zeropad3D_CP_2152_elements(402)); -- 
    -- CP-element group 403:  transition  input  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	391 
    -- CP-element group 403: successors 
    -- CP-element group 403:  members (5) 
      -- CP-element group 403: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Sample/word_access_start/word_0/$exit
      -- CP-element group 403: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Sample/word_access_start/$exit
      -- CP-element group 403: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Sample/$exit
      -- CP-element group 403: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_sample_completed_
      -- CP-element group 403: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Sample/word_access_start/word_0/ra
      -- 
    ra_6893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2954_load_0_ack_0, ack => zeropad3D_CP_2152_elements(403)); -- 
    -- CP-element group 404:  transition  input  output  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	391 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (12) 
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Update/LOAD_row_high_2954_Merge/$exit
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Update/LOAD_row_high_2954_Merge/$entry
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Update/word_access_complete/word_0/ca
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Update/word_access_complete/word_0/$exit
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Update/word_access_complete/$exit
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_update_completed_
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Update/$exit
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Update/LOAD_row_high_2954_Merge/merge_req
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/LOAD_row_high_2954_Update/LOAD_row_high_2954_Merge/merge_ack
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2958_sample_start_
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2958_Sample/$entry
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2958_Sample/rr
      -- 
    ca_6904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2954_load_0_ack_1, ack => zeropad3D_CP_2152_elements(404)); -- 
    rr_6917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(404), ack => type_cast_2958_inst_req_0); -- 
    -- CP-element group 405:  transition  input  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2958_sample_completed_
      -- CP-element group 405: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2958_Sample/$exit
      -- CP-element group 405: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2958_Sample/ra
      -- 
    ra_6918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2958_inst_ack_0, ack => zeropad3D_CP_2152_elements(405)); -- 
    -- CP-element group 406:  transition  input  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	391 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (3) 
      -- CP-element group 406: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2958_update_completed_
      -- CP-element group 406: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2958_Update/$exit
      -- CP-element group 406: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/type_cast_2958_Update/ca
      -- 
    ca_6923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2958_inst_ack_1, ack => zeropad3D_CP_2152_elements(406)); -- 
    -- CP-element group 407:  branch  join  transition  place  output  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	402 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407: 	409 
    -- CP-element group 407:  members (10) 
      -- CP-element group 407: 	 branch_block_stmt_714/if_stmt_2976__entry__
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975__exit__
      -- CP-element group 407: 	 branch_block_stmt_714/R_cmp828_2977_place
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2910_to_assign_stmt_2975/$exit
      -- CP-element group 407: 	 branch_block_stmt_714/if_stmt_2976_dead_link/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/if_stmt_2976_eval_test/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/if_stmt_2976_eval_test/$exit
      -- CP-element group 407: 	 branch_block_stmt_714/if_stmt_2976_eval_test/branch_req
      -- CP-element group 407: 	 branch_block_stmt_714/if_stmt_2976_if_link/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/if_stmt_2976_else_link/$entry
      -- 
    branch_req_6931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(407), ack => if_stmt_2976_branch_req_0); -- 
    zeropad3D_cp_element_group_407: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_407"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(402) & zeropad3D_CP_2152_elements(406);
      gj_zeropad3D_cp_element_group_407 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(407), clk => clk, reset => reset); --
    end block;
    -- CP-element group 408:  fork  transition  place  input  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	998 
    -- CP-element group 408: 	999 
    -- CP-element group 408: 	1001 
    -- CP-element group 408: 	1002 
    -- CP-element group 408:  members (20) 
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/type_cast_3012/SplitProtocol/Sample/$entry
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/type_cast_3012/SplitProtocol/Sample/rr
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/type_cast_3012/SplitProtocol/Update/$entry
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/type_cast_3012/SplitProtocol/Update/cr
      -- CP-element group 408: 	 branch_block_stmt_714/if_stmt_2976_if_link/$exit
      -- CP-element group 408: 	 branch_block_stmt_714/if_stmt_2976_if_link/if_choice_transition
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/$entry
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/$entry
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3008/SplitProtocol/Update/cr
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3008/SplitProtocol/Update/$entry
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3008/SplitProtocol/Sample/rr
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3008/SplitProtocol/Sample/$entry
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3008/SplitProtocol/$entry
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3008/$entry
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/$entry
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/$entry
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/$entry
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/type_cast_3012/SplitProtocol/$entry
      -- CP-element group 408: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/type_cast_3012/$entry
      -- 
    if_choice_transition_6936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2976_branch_ack_1, ack => zeropad3D_CP_2152_elements(408)); -- 
    rr_12630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(408), ack => type_cast_3012_inst_req_0); -- 
    cr_12635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(408), ack => type_cast_3012_inst_req_1); -- 
    cr_12612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(408), ack => type_cast_3008_inst_req_1); -- 
    rr_12607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(408), ack => type_cast_3008_inst_req_0); -- 
    -- CP-element group 409:  fork  transition  place  input  output  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	407 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	975 
    -- CP-element group 409: 	976 
    -- CP-element group 409: 	977 
    -- CP-element group 409: 	979 
    -- CP-element group 409: 	980 
    -- CP-element group 409:  members (22) 
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837
      -- CP-element group 409: 	 branch_block_stmt_714/if_stmt_2976_else_link/$exit
      -- CP-element group 409: 	 branch_block_stmt_714/if_stmt_2976_else_link/else_choice_transition
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_3001/SplitProtocol/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2983/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_3001/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2995/SplitProtocol/Update/cr
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2995/SplitProtocol/Update/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2995/SplitProtocol/Sample/rr
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2995/SplitProtocol/Sample/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2995/SplitProtocol/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2995/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_3001/SplitProtocol/Update/cr
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_3001/SplitProtocol/Update/$entry
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_3001/SplitProtocol/Sample/rr
      -- CP-element group 409: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_3001/SplitProtocol/Sample/$entry
      -- 
    else_choice_transition_6940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2976_branch_ack_0, ack => zeropad3D_CP_2152_elements(409)); -- 
    cr_12484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(409), ack => type_cast_2995_inst_req_1); -- 
    rr_12479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(409), ack => type_cast_2995_inst_req_0); -- 
    cr_12507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(409), ack => type_cast_3001_inst_req_1); -- 
    rr_12502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(409), ack => type_cast_3001_inst_req_0); -- 
    -- CP-element group 410:  transition  input  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	1007 
    -- CP-element group 410: successors 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3016_sample_completed_
      -- CP-element group 410: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3016_Sample/$exit
      -- CP-element group 410: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3016_Sample/ra
      -- 
    ra_6954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3016_inst_ack_0, ack => zeropad3D_CP_2152_elements(410)); -- 
    -- CP-element group 411:  transition  input  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	1007 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	424 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3016_update_completed_
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3016_Update/$exit
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3016_Update/ca
      -- 
    ca_6959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3016_inst_ack_1, ack => zeropad3D_CP_2152_elements(411)); -- 
    -- CP-element group 412:  transition  input  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	1007 
    -- CP-element group 412: successors 
    -- CP-element group 412:  members (5) 
      -- CP-element group 412: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_sample_completed_
      -- CP-element group 412: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Sample/$exit
      -- CP-element group 412: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Sample/word_access_start/$exit
      -- CP-element group 412: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Sample/word_access_start/word_0/$exit
      -- CP-element group 412: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Sample/word_access_start/word_0/ra
      -- 
    ra_6976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3025_load_0_ack_0, ack => zeropad3D_CP_2152_elements(412)); -- 
    -- CP-element group 413:  transition  input  output  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	1007 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	422 
    -- CP-element group 413:  members (12) 
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_update_completed_
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Update/$exit
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Update/word_access_complete/$exit
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Update/word_access_complete/word_0/$exit
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Update/word_access_complete/word_0/ca
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Update/LOAD_pad_3025_Merge/$entry
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Update/LOAD_pad_3025_Merge/$exit
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Update/LOAD_pad_3025_Merge/merge_req
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Update/LOAD_pad_3025_Merge/merge_ack
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3095_sample_start_
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3095_Sample/$entry
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3095_Sample/rr
      -- 
    ca_6987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3025_load_0_ack_1, ack => zeropad3D_CP_2152_elements(413)); -- 
    rr_7147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(413), ack => type_cast_3095_inst_req_0); -- 
    -- CP-element group 414:  transition  input  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	1007 
    -- CP-element group 414: successors 
    -- CP-element group 414:  members (5) 
      -- CP-element group 414: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_sample_completed_
      -- CP-element group 414: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Sample/$exit
      -- CP-element group 414: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Sample/word_access_start/$exit
      -- CP-element group 414: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Sample/word_access_start/word_0/$exit
      -- CP-element group 414: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Sample/word_access_start/word_0/ra
      -- 
    ra_7009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_3028_load_0_ack_0, ack => zeropad3D_CP_2152_elements(414)); -- 
    -- CP-element group 415:  transition  input  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	1007 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	420 
    -- CP-element group 415:  members (12) 
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_update_completed_
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Update/$exit
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Update/word_access_complete/$exit
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Update/word_access_complete/word_0/$exit
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Update/word_access_complete/word_0/ca
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Update/LOAD_depth_high_3028_Merge/$entry
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Update/LOAD_depth_high_3028_Merge/$exit
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Update/LOAD_depth_high_3028_Merge/merge_req
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Update/LOAD_depth_high_3028_Merge/merge_ack
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3056_sample_start_
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3056_Sample/$entry
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3056_Sample/rr
      -- 
    ca_7020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_3028_load_0_ack_1, ack => zeropad3D_CP_2152_elements(415)); -- 
    rr_7133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(415), ack => type_cast_3056_inst_req_0); -- 
    -- CP-element group 416:  transition  input  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	1007 
    -- CP-element group 416: successors 
    -- CP-element group 416:  members (5) 
      -- CP-element group 416: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_sample_completed_
      -- CP-element group 416: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Sample/$exit
      -- CP-element group 416: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Sample/word_access_start/$exit
      -- CP-element group 416: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Sample/word_access_start/word_0/$exit
      -- CP-element group 416: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Sample/word_access_start/word_0/ra
      -- 
    ra_7059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3040_load_0_ack_0, ack => zeropad3D_CP_2152_elements(416)); -- 
    -- CP-element group 417:  transition  input  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	1007 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	424 
    -- CP-element group 417:  members (9) 
      -- CP-element group 417: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_update_completed_
      -- CP-element group 417: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Update/$exit
      -- CP-element group 417: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Update/word_access_complete/$exit
      -- CP-element group 417: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Update/word_access_complete/word_0/$exit
      -- CP-element group 417: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Update/word_access_complete/word_0/ca
      -- CP-element group 417: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Update/ptr_deref_3040_Merge/$entry
      -- CP-element group 417: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Update/ptr_deref_3040_Merge/$exit
      -- CP-element group 417: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Update/ptr_deref_3040_Merge/merge_req
      -- CP-element group 417: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Update/ptr_deref_3040_Merge/merge_ack
      -- 
    ca_7070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3040_load_0_ack_1, ack => zeropad3D_CP_2152_elements(417)); -- 
    -- CP-element group 418:  transition  input  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	1007 
    -- CP-element group 418: successors 
    -- CP-element group 418:  members (5) 
      -- CP-element group 418: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_sample_completed_
      -- CP-element group 418: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Sample/$exit
      -- CP-element group 418: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Sample/word_access_start/$exit
      -- CP-element group 418: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Sample/word_access_start/word_0/$exit
      -- CP-element group 418: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Sample/word_access_start/word_0/ra
      -- 
    ra_7109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3052_load_0_ack_0, ack => zeropad3D_CP_2152_elements(418)); -- 
    -- CP-element group 419:  transition  input  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	1007 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	424 
    -- CP-element group 419:  members (9) 
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_update_completed_
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Update/$exit
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Update/word_access_complete/$exit
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Update/word_access_complete/word_0/$exit
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Update/word_access_complete/word_0/ca
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Update/ptr_deref_3052_Merge/$entry
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Update/ptr_deref_3052_Merge/$exit
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Update/ptr_deref_3052_Merge/merge_req
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Update/ptr_deref_3052_Merge/merge_ack
      -- 
    ca_7120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3052_load_0_ack_1, ack => zeropad3D_CP_2152_elements(419)); -- 
    -- CP-element group 420:  transition  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	415 
    -- CP-element group 420: successors 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3056_sample_completed_
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3056_Sample/$exit
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3056_Sample/ra
      -- 
    ra_7134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3056_inst_ack_0, ack => zeropad3D_CP_2152_elements(420)); -- 
    -- CP-element group 421:  transition  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	1007 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	424 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3056_update_completed_
      -- CP-element group 421: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3056_Update/$exit
      -- CP-element group 421: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3056_Update/ca
      -- 
    ca_7139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3056_inst_ack_1, ack => zeropad3D_CP_2152_elements(421)); -- 
    -- CP-element group 422:  transition  input  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	413 
    -- CP-element group 422: successors 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3095_sample_completed_
      -- CP-element group 422: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3095_Sample/$exit
      -- CP-element group 422: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3095_Sample/ra
      -- 
    ra_7148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3095_inst_ack_0, ack => zeropad3D_CP_2152_elements(422)); -- 
    -- CP-element group 423:  transition  input  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	1007 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3095_update_completed_
      -- CP-element group 423: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3095_Update/$exit
      -- CP-element group 423: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3095_Update/ca
      -- 
    ca_7153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3095_inst_ack_1, ack => zeropad3D_CP_2152_elements(423)); -- 
    -- CP-element group 424:  join  fork  transition  place  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	411 
    -- CP-element group 424: 	417 
    -- CP-element group 424: 	419 
    -- CP-element group 424: 	421 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	1018 
    -- CP-element group 424: 	1019 
    -- CP-element group 424: 	1020 
    -- CP-element group 424: 	1022 
    -- CP-element group 424:  members (16) 
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137__exit__
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/$exit
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3153/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3152/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3140/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3152/SplitProtocol/Update/cr
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3152/SplitProtocol/Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3152/SplitProtocol/Sample/rr
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3152/SplitProtocol/Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3152/SplitProtocol/$entry
      -- 
    cr_12747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => type_cast_3152_inst_req_1); -- 
    rr_12742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => type_cast_3152_inst_req_0); -- 
    zeropad3D_cp_element_group_424: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_424"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(411) & zeropad3D_CP_2152_elements(417) & zeropad3D_CP_2152_elements(419) & zeropad3D_CP_2152_elements(421) & zeropad3D_CP_2152_elements(423);
      gj_zeropad3D_cp_element_group_424 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(424), clk => clk, reset => reset); --
    end block;
    -- CP-element group 425:  transition  input  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	1028 
    -- CP-element group 425: successors 
    -- CP-element group 425:  members (3) 
      -- CP-element group 425: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/type_cast_3164_sample_completed_
      -- CP-element group 425: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/type_cast_3164_Sample/$exit
      -- CP-element group 425: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/type_cast_3164_Sample/ra
      -- 
    ra_7165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3164_inst_ack_0, ack => zeropad3D_CP_2152_elements(425)); -- 
    -- CP-element group 426:  branch  transition  place  input  output  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	1028 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426: 	428 
    -- CP-element group 426:  members (13) 
      -- CP-element group 426: 	 branch_block_stmt_714/if_stmt_3173__entry__
      -- CP-element group 426: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172__exit__
      -- CP-element group 426: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/$exit
      -- CP-element group 426: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/type_cast_3164_update_completed_
      -- CP-element group 426: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/type_cast_3164_Update/$exit
      -- CP-element group 426: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/type_cast_3164_Update/ca
      -- CP-element group 426: 	 branch_block_stmt_714/if_stmt_3173_dead_link/$entry
      -- CP-element group 426: 	 branch_block_stmt_714/if_stmt_3173_eval_test/$entry
      -- CP-element group 426: 	 branch_block_stmt_714/if_stmt_3173_eval_test/$exit
      -- CP-element group 426: 	 branch_block_stmt_714/if_stmt_3173_eval_test/branch_req
      -- CP-element group 426: 	 branch_block_stmt_714/R_cmp903_3174_place
      -- CP-element group 426: 	 branch_block_stmt_714/if_stmt_3173_if_link/$entry
      -- CP-element group 426: 	 branch_block_stmt_714/if_stmt_3173_else_link/$entry
      -- 
    ca_7170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3164_inst_ack_1, ack => zeropad3D_CP_2152_elements(426)); -- 
    branch_req_7178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(426), ack => if_stmt_3173_branch_req_0); -- 
    -- CP-element group 427:  transition  place  input  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	1029 
    -- CP-element group 427:  members (5) 
      -- CP-element group 427: 	 branch_block_stmt_714/if_stmt_3173_if_link/$exit
      -- CP-element group 427: 	 branch_block_stmt_714/if_stmt_3173_if_link/if_choice_transition
      -- CP-element group 427: 	 branch_block_stmt_714/whilex_xbody898_ifx_xthen935
      -- CP-element group 427: 	 branch_block_stmt_714/whilex_xbody898_ifx_xthen935_PhiReq/$entry
      -- CP-element group 427: 	 branch_block_stmt_714/whilex_xbody898_ifx_xthen935_PhiReq/$exit
      -- 
    if_choice_transition_7183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3173_branch_ack_1, ack => zeropad3D_CP_2152_elements(427)); -- 
    -- CP-element group 428:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	426 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	429 
    -- CP-element group 428: 	430 
    -- CP-element group 428: 	432 
    -- CP-element group 428:  members (27) 
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210__entry__
      -- CP-element group 428: 	 branch_block_stmt_714/merge_stmt_3179__exit__
      -- CP-element group 428: 	 branch_block_stmt_714/if_stmt_3173_else_link/$exit
      -- CP-element group 428: 	 branch_block_stmt_714/if_stmt_3173_else_link/else_choice_transition
      -- CP-element group 428: 	 branch_block_stmt_714/whilex_xbody898_lorx_xlhsx_xfalse905
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/$entry
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_sample_start_
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_update_start_
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_word_address_calculated
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_root_address_calculated
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Sample/$entry
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Sample/word_access_start/$entry
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Sample/word_access_start/word_0/$entry
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Sample/word_access_start/word_0/rr
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Update/$entry
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Update/word_access_complete/$entry
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Update/word_access_complete/word_0/$entry
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Update/word_access_complete/word_0/cr
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/type_cast_3185_update_start_
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/type_cast_3185_Update/$entry
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/type_cast_3185_Update/cr
      -- CP-element group 428: 	 branch_block_stmt_714/merge_stmt_3179_PhiAck/$entry
      -- CP-element group 428: 	 branch_block_stmt_714/merge_stmt_3179_PhiReqMerge
      -- CP-element group 428: 	 branch_block_stmt_714/whilex_xbody898_lorx_xlhsx_xfalse905_PhiReq/$exit
      -- CP-element group 428: 	 branch_block_stmt_714/whilex_xbody898_lorx_xlhsx_xfalse905_PhiReq/$entry
      -- CP-element group 428: 	 branch_block_stmt_714/merge_stmt_3179_PhiAck/dummy
      -- CP-element group 428: 	 branch_block_stmt_714/merge_stmt_3179_PhiAck/$exit
      -- 
    else_choice_transition_7187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3173_branch_ack_0, ack => zeropad3D_CP_2152_elements(428)); -- 
    rr_7208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(428), ack => LOAD_row_high_3181_load_0_req_0); -- 
    cr_7219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(428), ack => LOAD_row_high_3181_load_0_req_1); -- 
    cr_7238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(428), ack => type_cast_3185_inst_req_1); -- 
    -- CP-element group 429:  transition  input  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	428 
    -- CP-element group 429: successors 
    -- CP-element group 429:  members (5) 
      -- CP-element group 429: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_sample_completed_
      -- CP-element group 429: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Sample/$exit
      -- CP-element group 429: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Sample/word_access_start/$exit
      -- CP-element group 429: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Sample/word_access_start/word_0/$exit
      -- CP-element group 429: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Sample/word_access_start/word_0/ra
      -- 
    ra_7209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3181_load_0_ack_0, ack => zeropad3D_CP_2152_elements(429)); -- 
    -- CP-element group 430:  transition  input  output  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	428 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	431 
    -- CP-element group 430:  members (12) 
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_update_completed_
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Update/$exit
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Update/word_access_complete/$exit
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Update/word_access_complete/word_0/$exit
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Update/word_access_complete/word_0/ca
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Update/LOAD_row_high_3181_Merge/$entry
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Update/LOAD_row_high_3181_Merge/$exit
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Update/LOAD_row_high_3181_Merge/merge_req
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/LOAD_row_high_3181_Update/LOAD_row_high_3181_Merge/merge_ack
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/type_cast_3185_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/type_cast_3185_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/type_cast_3185_Sample/rr
      -- 
    ca_7220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3181_load_0_ack_1, ack => zeropad3D_CP_2152_elements(430)); -- 
    rr_7233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(430), ack => type_cast_3185_inst_req_0); -- 
    -- CP-element group 431:  transition  input  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	430 
    -- CP-element group 431: successors 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/type_cast_3185_sample_completed_
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/type_cast_3185_Sample/$exit
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/type_cast_3185_Sample/ra
      -- 
    ra_7234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3185_inst_ack_0, ack => zeropad3D_CP_2152_elements(431)); -- 
    -- CP-element group 432:  branch  transition  place  input  output  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	428 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	433 
    -- CP-element group 432: 	434 
    -- CP-element group 432:  members (13) 
      -- CP-element group 432: 	 branch_block_stmt_714/if_stmt_3211__entry__
      -- CP-element group 432: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210__exit__
      -- CP-element group 432: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/$exit
      -- CP-element group 432: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/type_cast_3185_update_completed_
      -- CP-element group 432: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/type_cast_3185_Update/$exit
      -- CP-element group 432: 	 branch_block_stmt_714/assign_stmt_3182_to_assign_stmt_3210/type_cast_3185_Update/ca
      -- CP-element group 432: 	 branch_block_stmt_714/if_stmt_3211_dead_link/$entry
      -- CP-element group 432: 	 branch_block_stmt_714/if_stmt_3211_eval_test/$entry
      -- CP-element group 432: 	 branch_block_stmt_714/if_stmt_3211_eval_test/$exit
      -- CP-element group 432: 	 branch_block_stmt_714/if_stmt_3211_eval_test/branch_req
      -- CP-element group 432: 	 branch_block_stmt_714/R_cmp915_3212_place
      -- CP-element group 432: 	 branch_block_stmt_714/if_stmt_3211_if_link/$entry
      -- CP-element group 432: 	 branch_block_stmt_714/if_stmt_3211_else_link/$entry
      -- 
    ca_7239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3185_inst_ack_1, ack => zeropad3D_CP_2152_elements(432)); -- 
    branch_req_7247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(432), ack => if_stmt_3211_branch_req_0); -- 
    -- CP-element group 433:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	432 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	435 
    -- CP-element group 433: 	436 
    -- CP-element group 433:  members (18) 
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229__entry__
      -- CP-element group 433: 	 branch_block_stmt_714/merge_stmt_3217__exit__
      -- CP-element group 433: 	 branch_block_stmt_714/if_stmt_3211_if_link/$exit
      -- CP-element group 433: 	 branch_block_stmt_714/if_stmt_3211_if_link/if_choice_transition
      -- CP-element group 433: 	 branch_block_stmt_714/lorx_xlhsx_xfalse905_lorx_xlhsx_xfalse917
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/$entry
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/type_cast_3221_sample_start_
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/type_cast_3221_update_start_
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/type_cast_3221_Sample/$entry
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/type_cast_3221_Sample/rr
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/type_cast_3221_Update/$entry
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/type_cast_3221_Update/cr
      -- CP-element group 433: 	 branch_block_stmt_714/merge_stmt_3217_PhiReqMerge
      -- CP-element group 433: 	 branch_block_stmt_714/lorx_xlhsx_xfalse905_lorx_xlhsx_xfalse917_PhiReq/$exit
      -- CP-element group 433: 	 branch_block_stmt_714/lorx_xlhsx_xfalse905_lorx_xlhsx_xfalse917_PhiReq/$entry
      -- CP-element group 433: 	 branch_block_stmt_714/merge_stmt_3217_PhiAck/$entry
      -- CP-element group 433: 	 branch_block_stmt_714/merge_stmt_3217_PhiAck/$exit
      -- CP-element group 433: 	 branch_block_stmt_714/merge_stmt_3217_PhiAck/dummy
      -- 
    if_choice_transition_7252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3211_branch_ack_1, ack => zeropad3D_CP_2152_elements(433)); -- 
    rr_7269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(433), ack => type_cast_3221_inst_req_0); -- 
    cr_7274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(433), ack => type_cast_3221_inst_req_1); -- 
    -- CP-element group 434:  transition  place  input  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	432 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	1029 
    -- CP-element group 434:  members (5) 
      -- CP-element group 434: 	 branch_block_stmt_714/if_stmt_3211_else_link/$exit
      -- CP-element group 434: 	 branch_block_stmt_714/if_stmt_3211_else_link/else_choice_transition
      -- CP-element group 434: 	 branch_block_stmt_714/lorx_xlhsx_xfalse905_ifx_xthen935
      -- CP-element group 434: 	 branch_block_stmt_714/lorx_xlhsx_xfalse905_ifx_xthen935_PhiReq/$entry
      -- CP-element group 434: 	 branch_block_stmt_714/lorx_xlhsx_xfalse905_ifx_xthen935_PhiReq/$exit
      -- 
    else_choice_transition_7256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3211_branch_ack_0, ack => zeropad3D_CP_2152_elements(434)); -- 
    -- CP-element group 435:  transition  input  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	433 
    -- CP-element group 435: successors 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/type_cast_3221_sample_completed_
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/type_cast_3221_Sample/$exit
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/type_cast_3221_Sample/ra
      -- 
    ra_7270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3221_inst_ack_0, ack => zeropad3D_CP_2152_elements(435)); -- 
    -- CP-element group 436:  branch  transition  place  input  output  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	433 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	437 
    -- CP-element group 436: 	438 
    -- CP-element group 436:  members (13) 
      -- CP-element group 436: 	 branch_block_stmt_714/if_stmt_3230__entry__
      -- CP-element group 436: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229__exit__
      -- CP-element group 436: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/$exit
      -- CP-element group 436: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/type_cast_3221_update_completed_
      -- CP-element group 436: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/type_cast_3221_Update/$exit
      -- CP-element group 436: 	 branch_block_stmt_714/assign_stmt_3222_to_assign_stmt_3229/type_cast_3221_Update/ca
      -- CP-element group 436: 	 branch_block_stmt_714/if_stmt_3230_dead_link/$entry
      -- CP-element group 436: 	 branch_block_stmt_714/if_stmt_3230_eval_test/$entry
      -- CP-element group 436: 	 branch_block_stmt_714/if_stmt_3230_eval_test/$exit
      -- CP-element group 436: 	 branch_block_stmt_714/if_stmt_3230_eval_test/branch_req
      -- CP-element group 436: 	 branch_block_stmt_714/R_cmp922_3231_place
      -- CP-element group 436: 	 branch_block_stmt_714/if_stmt_3230_if_link/$entry
      -- CP-element group 436: 	 branch_block_stmt_714/if_stmt_3230_else_link/$entry
      -- 
    ca_7275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3221_inst_ack_1, ack => zeropad3D_CP_2152_elements(436)); -- 
    branch_req_7283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(436), ack => if_stmt_3230_branch_req_0); -- 
    -- CP-element group 437:  transition  place  input  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	436 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	1029 
    -- CP-element group 437:  members (5) 
      -- CP-element group 437: 	 branch_block_stmt_714/if_stmt_3230_if_link/$exit
      -- CP-element group 437: 	 branch_block_stmt_714/if_stmt_3230_if_link/if_choice_transition
      -- CP-element group 437: 	 branch_block_stmt_714/lorx_xlhsx_xfalse917_ifx_xthen935
      -- CP-element group 437: 	 branch_block_stmt_714/lorx_xlhsx_xfalse917_ifx_xthen935_PhiReq/$entry
      -- CP-element group 437: 	 branch_block_stmt_714/lorx_xlhsx_xfalse917_ifx_xthen935_PhiReq/$exit
      -- 
    if_choice_transition_7288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3230_branch_ack_1, ack => zeropad3D_CP_2152_elements(437)); -- 
    -- CP-element group 438:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	436 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	439 
    -- CP-element group 438: 	440 
    -- CP-element group 438: 	442 
    -- CP-element group 438:  members (27) 
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261__entry__
      -- CP-element group 438: 	 branch_block_stmt_714/merge_stmt_3236__exit__
      -- CP-element group 438: 	 branch_block_stmt_714/if_stmt_3230_else_link/$exit
      -- CP-element group 438: 	 branch_block_stmt_714/if_stmt_3230_else_link/else_choice_transition
      -- CP-element group 438: 	 branch_block_stmt_714/lorx_xlhsx_xfalse917_lorx_xlhsx_xfalse924
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/$entry
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_sample_start_
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_update_start_
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_word_address_calculated
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_root_address_calculated
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Sample/$entry
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Sample/word_access_start/$entry
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Sample/word_access_start/word_0/$entry
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Sample/word_access_start/word_0/rr
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Update/word_access_complete/$entry
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Update/word_access_complete/word_0/$entry
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Update/word_access_complete/word_0/cr
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/type_cast_3242_update_start_
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/type_cast_3242_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/type_cast_3242_Update/cr
      -- CP-element group 438: 	 branch_block_stmt_714/lorx_xlhsx_xfalse917_lorx_xlhsx_xfalse924_PhiReq/$entry
      -- CP-element group 438: 	 branch_block_stmt_714/lorx_xlhsx_xfalse917_lorx_xlhsx_xfalse924_PhiReq/$exit
      -- CP-element group 438: 	 branch_block_stmt_714/merge_stmt_3236_PhiReqMerge
      -- CP-element group 438: 	 branch_block_stmt_714/merge_stmt_3236_PhiAck/$entry
      -- CP-element group 438: 	 branch_block_stmt_714/merge_stmt_3236_PhiAck/$exit
      -- CP-element group 438: 	 branch_block_stmt_714/merge_stmt_3236_PhiAck/dummy
      -- 
    else_choice_transition_7292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3230_branch_ack_0, ack => zeropad3D_CP_2152_elements(438)); -- 
    rr_7313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(438), ack => LOAD_col_high_3238_load_0_req_0); -- 
    cr_7324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(438), ack => LOAD_col_high_3238_load_0_req_1); -- 
    cr_7343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(438), ack => type_cast_3242_inst_req_1); -- 
    -- CP-element group 439:  transition  input  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	438 
    -- CP-element group 439: successors 
    -- CP-element group 439:  members (5) 
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_sample_completed_
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Sample/$exit
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Sample/word_access_start/$exit
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Sample/word_access_start/word_0/$exit
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Sample/word_access_start/word_0/ra
      -- 
    ra_7314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3238_load_0_ack_0, ack => zeropad3D_CP_2152_elements(439)); -- 
    -- CP-element group 440:  transition  input  output  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	438 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	441 
    -- CP-element group 440:  members (12) 
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_update_completed_
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Update/$exit
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Update/word_access_complete/$exit
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Update/word_access_complete/word_0/$exit
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Update/word_access_complete/word_0/ca
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Update/LOAD_col_high_3238_Merge/$entry
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Update/LOAD_col_high_3238_Merge/$exit
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Update/LOAD_col_high_3238_Merge/merge_req
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/LOAD_col_high_3238_Update/LOAD_col_high_3238_Merge/merge_ack
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/type_cast_3242_sample_start_
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/type_cast_3242_Sample/$entry
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/type_cast_3242_Sample/rr
      -- 
    ca_7325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3238_load_0_ack_1, ack => zeropad3D_CP_2152_elements(440)); -- 
    rr_7338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(440), ack => type_cast_3242_inst_req_0); -- 
    -- CP-element group 441:  transition  input  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	440 
    -- CP-element group 441: successors 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/type_cast_3242_sample_completed_
      -- CP-element group 441: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/type_cast_3242_Sample/$exit
      -- CP-element group 441: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/type_cast_3242_Sample/ra
      -- 
    ra_7339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3242_inst_ack_0, ack => zeropad3D_CP_2152_elements(441)); -- 
    -- CP-element group 442:  branch  transition  place  input  output  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	438 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	443 
    -- CP-element group 442: 	444 
    -- CP-element group 442:  members (13) 
      -- CP-element group 442: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261__exit__
      -- CP-element group 442: 	 branch_block_stmt_714/if_stmt_3262__entry__
      -- CP-element group 442: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/$exit
      -- CP-element group 442: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/type_cast_3242_update_completed_
      -- CP-element group 442: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/type_cast_3242_Update/$exit
      -- CP-element group 442: 	 branch_block_stmt_714/assign_stmt_3239_to_assign_stmt_3261/type_cast_3242_Update/ca
      -- CP-element group 442: 	 branch_block_stmt_714/if_stmt_3262_dead_link/$entry
      -- CP-element group 442: 	 branch_block_stmt_714/if_stmt_3262_eval_test/$entry
      -- CP-element group 442: 	 branch_block_stmt_714/if_stmt_3262_eval_test/$exit
      -- CP-element group 442: 	 branch_block_stmt_714/if_stmt_3262_eval_test/branch_req
      -- CP-element group 442: 	 branch_block_stmt_714/R_cmp933_3263_place
      -- CP-element group 442: 	 branch_block_stmt_714/if_stmt_3262_if_link/$entry
      -- CP-element group 442: 	 branch_block_stmt_714/if_stmt_3262_else_link/$entry
      -- 
    ca_7344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3242_inst_ack_1, ack => zeropad3D_CP_2152_elements(442)); -- 
    branch_req_7352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(442), ack => if_stmt_3262_branch_req_0); -- 
    -- CP-element group 443:  fork  transition  place  input  output  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	442 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	459 
    -- CP-element group 443: 	460 
    -- CP-element group 443: 	462 
    -- CP-element group 443: 	464 
    -- CP-element group 443: 	466 
    -- CP-element group 443: 	468 
    -- CP-element group 443: 	470 
    -- CP-element group 443: 	472 
    -- CP-element group 443: 	474 
    -- CP-element group 443: 	477 
    -- CP-element group 443:  members (46) 
      -- CP-element group 443: 	 branch_block_stmt_714/merge_stmt_3326__exit__
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431__entry__
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_update_start_
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Update/word_access_complete/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3426_complete/req
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3426_complete/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Update/word_access_complete/word_0/cr
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Update/word_access_complete/word_0/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/if_stmt_3262_if_link/$exit
      -- CP-element group 443: 	 branch_block_stmt_714/if_stmt_3262_if_link/if_choice_transition
      -- CP-element group 443: 	 branch_block_stmt_714/lorx_xlhsx_xfalse924_ifx_xelse956
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3330_sample_start_
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3330_update_start_
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3330_Sample/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3330_Sample/rr
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3330_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3330_Update/cr
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3394_update_start_
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3394_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3394_Update/cr
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3401_update_start_
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_final_index_sum_regn_update_start
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_final_index_sum_regn_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_final_index_sum_regn_Update/req
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3401_complete/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3401_complete/req
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_update_start_
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Update/word_access_complete/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Update/word_access_complete/word_0/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Update/word_access_complete/word_0/cr
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3419_update_start_
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3419_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3419_Update/cr
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3426_update_start_
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_final_index_sum_regn_update_start
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_final_index_sum_regn_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_final_index_sum_regn_Update/req
      -- CP-element group 443: 	 branch_block_stmt_714/lorx_xlhsx_xfalse924_ifx_xelse956_PhiReq/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/lorx_xlhsx_xfalse924_ifx_xelse956_PhiReq/$exit
      -- CP-element group 443: 	 branch_block_stmt_714/merge_stmt_3326_PhiReqMerge
      -- CP-element group 443: 	 branch_block_stmt_714/merge_stmt_3326_PhiAck/$entry
      -- CP-element group 443: 	 branch_block_stmt_714/merge_stmt_3326_PhiAck/$exit
      -- CP-element group 443: 	 branch_block_stmt_714/merge_stmt_3326_PhiAck/dummy
      -- 
    if_choice_transition_7357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3262_branch_ack_1, ack => zeropad3D_CP_2152_elements(443)); -- 
    req_7690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(443), ack => addr_of_3426_final_reg_req_1); -- 
    cr_7740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(443), ack => ptr_deref_3429_store_0_req_1); -- 
    rr_7515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(443), ack => type_cast_3330_inst_req_0); -- 
    cr_7520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(443), ack => type_cast_3330_inst_req_1); -- 
    cr_7534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(443), ack => type_cast_3394_inst_req_1); -- 
    req_7565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(443), ack => array_obj_ref_3400_index_offset_req_1); -- 
    req_7580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(443), ack => addr_of_3401_final_reg_req_1); -- 
    cr_7625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(443), ack => ptr_deref_3405_load_0_req_1); -- 
    cr_7644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(443), ack => type_cast_3419_inst_req_1); -- 
    req_7675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(443), ack => array_obj_ref_3425_index_offset_req_1); -- 
    -- CP-element group 444:  transition  place  input  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	442 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	1029 
    -- CP-element group 444:  members (5) 
      -- CP-element group 444: 	 branch_block_stmt_714/if_stmt_3262_else_link/$exit
      -- CP-element group 444: 	 branch_block_stmt_714/if_stmt_3262_else_link/else_choice_transition
      -- CP-element group 444: 	 branch_block_stmt_714/lorx_xlhsx_xfalse924_ifx_xthen935
      -- CP-element group 444: 	 branch_block_stmt_714/lorx_xlhsx_xfalse924_ifx_xthen935_PhiReq/$entry
      -- CP-element group 444: 	 branch_block_stmt_714/lorx_xlhsx_xfalse924_ifx_xthen935_PhiReq/$exit
      -- 
    else_choice_transition_7361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3262_branch_ack_0, ack => zeropad3D_CP_2152_elements(444)); -- 
    -- CP-element group 445:  transition  input  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	1029 
    -- CP-element group 445: successors 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3272_sample_completed_
      -- CP-element group 445: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3272_Sample/$exit
      -- CP-element group 445: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3272_Sample/ra
      -- 
    ra_7375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3272_inst_ack_0, ack => zeropad3D_CP_2152_elements(445)); -- 
    -- CP-element group 446:  transition  input  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	1029 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	449 
    -- CP-element group 446:  members (3) 
      -- CP-element group 446: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3272_update_completed_
      -- CP-element group 446: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3272_Update/$exit
      -- CP-element group 446: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3272_Update/ca
      -- 
    ca_7380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3272_inst_ack_1, ack => zeropad3D_CP_2152_elements(446)); -- 
    -- CP-element group 447:  transition  input  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	1029 
    -- CP-element group 447: successors 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3277_sample_completed_
      -- CP-element group 447: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3277_Sample/$exit
      -- CP-element group 447: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3277_Sample/ra
      -- 
    ra_7389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3277_inst_ack_0, ack => zeropad3D_CP_2152_elements(447)); -- 
    -- CP-element group 448:  transition  input  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	1029 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (3) 
      -- CP-element group 448: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3277_update_completed_
      -- CP-element group 448: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3277_Update/$exit
      -- CP-element group 448: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3277_Update/ca
      -- 
    ca_7394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3277_inst_ack_1, ack => zeropad3D_CP_2152_elements(448)); -- 
    -- CP-element group 449:  join  transition  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	446 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	450 
    -- CP-element group 449:  members (3) 
      -- CP-element group 449: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3311_sample_start_
      -- CP-element group 449: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3311_Sample/$entry
      -- CP-element group 449: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3311_Sample/rr
      -- 
    rr_7402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(449), ack => type_cast_3311_inst_req_0); -- 
    zeropad3D_cp_element_group_449: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_449"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(446) & zeropad3D_CP_2152_elements(448);
      gj_zeropad3D_cp_element_group_449 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 450:  transition  input  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	449 
    -- CP-element group 450: successors 
    -- CP-element group 450:  members (3) 
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3311_sample_completed_
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3311_Sample/$exit
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3311_Sample/ra
      -- 
    ra_7403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3311_inst_ack_0, ack => zeropad3D_CP_2152_elements(450)); -- 
    -- CP-element group 451:  transition  input  output  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	1029 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	452 
    -- CP-element group 451:  members (16) 
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3311_update_completed_
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3311_Update/$exit
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3311_Update/ca
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_index_resized_1
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_index_scaled_1
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_index_computed_1
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_index_resize_1/$entry
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_index_resize_1/$exit
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_index_resize_1/index_resize_req
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_index_resize_1/index_resize_ack
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_index_scale_1/$entry
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_index_scale_1/$exit
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_index_scale_1/scale_rename_req
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_index_scale_1/scale_rename_ack
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_final_index_sum_regn_Sample/$entry
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_final_index_sum_regn_Sample/req
      -- 
    ca_7408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3311_inst_ack_1, ack => zeropad3D_CP_2152_elements(451)); -- 
    req_7433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(451), ack => array_obj_ref_3317_index_offset_req_0); -- 
    -- CP-element group 452:  transition  input  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	451 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	458 
    -- CP-element group 452:  members (3) 
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_final_index_sum_regn_sample_complete
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_final_index_sum_regn_Sample/$exit
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_final_index_sum_regn_Sample/ack
      -- 
    ack_7434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3317_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(452)); -- 
    -- CP-element group 453:  transition  input  output  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	1029 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	454 
    -- CP-element group 453:  members (11) 
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/addr_of_3318_sample_start_
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_root_address_calculated
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_offset_calculated
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_final_index_sum_regn_Update/$exit
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_final_index_sum_regn_Update/ack
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_base_plus_offset/$entry
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_base_plus_offset/$exit
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_base_plus_offset/sum_rename_req
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_base_plus_offset/sum_rename_ack
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/addr_of_3318_request/$entry
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/addr_of_3318_request/req
      -- 
    ack_7439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3317_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(453)); -- 
    req_7448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(453), ack => addr_of_3318_final_reg_req_0); -- 
    -- CP-element group 454:  transition  input  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	453 
    -- CP-element group 454: successors 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/addr_of_3318_sample_completed_
      -- CP-element group 454: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/addr_of_3318_request/$exit
      -- CP-element group 454: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/addr_of_3318_request/ack
      -- 
    ack_7449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3318_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(454)); -- 
    -- CP-element group 455:  join  fork  transition  input  output  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	1029 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455:  members (28) 
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/addr_of_3318_update_completed_
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/addr_of_3318_complete/$exit
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/addr_of_3318_complete/ack
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_sample_start_
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_base_address_calculated
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_word_address_calculated
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_root_address_calculated
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_base_address_resized
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_base_addr_resize/$entry
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_base_addr_resize/$exit
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_base_addr_resize/base_resize_req
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_base_addr_resize/base_resize_ack
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_base_plus_offset/$entry
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_base_plus_offset/$exit
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_base_plus_offset/sum_rename_req
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_base_plus_offset/sum_rename_ack
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_word_addrgen/$entry
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_word_addrgen/$exit
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_word_addrgen/root_register_req
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_word_addrgen/root_register_ack
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Sample/$entry
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Sample/ptr_deref_3321_Split/$entry
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Sample/ptr_deref_3321_Split/$exit
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Sample/ptr_deref_3321_Split/split_req
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Sample/ptr_deref_3321_Split/split_ack
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Sample/word_access_start/$entry
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Sample/word_access_start/word_0/$entry
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Sample/word_access_start/word_0/rr
      -- 
    ack_7454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3318_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(455)); -- 
    rr_7492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(455), ack => ptr_deref_3321_store_0_req_0); -- 
    -- CP-element group 456:  transition  input  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	455 
    -- CP-element group 456: successors 
    -- CP-element group 456:  members (5) 
      -- CP-element group 456: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_sample_completed_
      -- CP-element group 456: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Sample/$exit
      -- CP-element group 456: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Sample/word_access_start/$exit
      -- CP-element group 456: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Sample/word_access_start/word_0/$exit
      -- CP-element group 456: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Sample/word_access_start/word_0/ra
      -- 
    ra_7493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3321_store_0_ack_0, ack => zeropad3D_CP_2152_elements(456)); -- 
    -- CP-element group 457:  transition  input  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	1029 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	458 
    -- CP-element group 457:  members (5) 
      -- CP-element group 457: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_update_completed_
      -- CP-element group 457: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Update/$exit
      -- CP-element group 457: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Update/word_access_complete/$exit
      -- CP-element group 457: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Update/word_access_complete/word_0/$exit
      -- CP-element group 457: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Update/word_access_complete/word_0/ca
      -- 
    ca_7504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 457_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3321_store_0_ack_1, ack => zeropad3D_CP_2152_elements(457)); -- 
    -- CP-element group 458:  join  transition  place  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	452 
    -- CP-element group 458: 	457 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	1030 
    -- CP-element group 458:  members (5) 
      -- CP-element group 458: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324__exit__
      -- CP-element group 458: 	 branch_block_stmt_714/ifx_xthen935_ifx_xend1004
      -- CP-element group 458: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/$exit
      -- CP-element group 458: 	 branch_block_stmt_714/ifx_xthen935_ifx_xend1004_PhiReq/$entry
      -- CP-element group 458: 	 branch_block_stmt_714/ifx_xthen935_ifx_xend1004_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_458: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_458"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(452) & zeropad3D_CP_2152_elements(457);
      gj_zeropad3D_cp_element_group_458 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(458), clk => clk, reset => reset); --
    end block;
    -- CP-element group 459:  transition  input  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	443 
    -- CP-element group 459: successors 
    -- CP-element group 459:  members (3) 
      -- CP-element group 459: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3330_sample_completed_
      -- CP-element group 459: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3330_Sample/$exit
      -- CP-element group 459: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3330_Sample/ra
      -- 
    ra_7516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3330_inst_ack_0, ack => zeropad3D_CP_2152_elements(459)); -- 
    -- CP-element group 460:  fork  transition  input  output  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	443 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	461 
    -- CP-element group 460: 	469 
    -- CP-element group 460:  members (9) 
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3330_update_completed_
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3330_Update/$exit
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3330_Update/ca
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3394_sample_start_
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3394_Sample/$entry
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3394_Sample/rr
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3419_sample_start_
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3419_Sample/$entry
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3419_Sample/rr
      -- 
    ca_7521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3330_inst_ack_1, ack => zeropad3D_CP_2152_elements(460)); -- 
    rr_7529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(460), ack => type_cast_3394_inst_req_0); -- 
    rr_7639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(460), ack => type_cast_3419_inst_req_0); -- 
    -- CP-element group 461:  transition  input  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	460 
    -- CP-element group 461: successors 
    -- CP-element group 461:  members (3) 
      -- CP-element group 461: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3394_sample_completed_
      -- CP-element group 461: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3394_Sample/$exit
      -- CP-element group 461: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3394_Sample/ra
      -- 
    ra_7530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3394_inst_ack_0, ack => zeropad3D_CP_2152_elements(461)); -- 
    -- CP-element group 462:  transition  input  output  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	443 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	463 
    -- CP-element group 462:  members (16) 
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3394_update_completed_
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3394_Update/$exit
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3394_Update/ca
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_index_resized_1
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_index_scaled_1
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_index_computed_1
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_index_resize_1/$entry
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_index_resize_1/$exit
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_index_resize_1/index_resize_req
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_index_resize_1/index_resize_ack
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_index_scale_1/$entry
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_index_scale_1/$exit
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_index_scale_1/scale_rename_req
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_index_scale_1/scale_rename_ack
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_final_index_sum_regn_Sample/$entry
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_final_index_sum_regn_Sample/req
      -- 
    ca_7535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3394_inst_ack_1, ack => zeropad3D_CP_2152_elements(462)); -- 
    req_7560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(462), ack => array_obj_ref_3400_index_offset_req_0); -- 
    -- CP-element group 463:  transition  input  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	462 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	478 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_final_index_sum_regn_sample_complete
      -- CP-element group 463: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_final_index_sum_regn_Sample/$exit
      -- CP-element group 463: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_final_index_sum_regn_Sample/ack
      -- 
    ack_7561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3400_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(463)); -- 
    -- CP-element group 464:  transition  input  output  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	443 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	465 
    -- CP-element group 464:  members (11) 
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3401_sample_start_
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_root_address_calculated
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_offset_calculated
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_final_index_sum_regn_Update/$exit
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_final_index_sum_regn_Update/ack
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_base_plus_offset/$entry
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_base_plus_offset/$exit
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_base_plus_offset/sum_rename_req
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3400_base_plus_offset/sum_rename_ack
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3401_request/$entry
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3401_request/req
      -- 
    ack_7566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3400_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(464)); -- 
    req_7575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(464), ack => addr_of_3401_final_reg_req_0); -- 
    -- CP-element group 465:  transition  input  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	464 
    -- CP-element group 465: successors 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3401_sample_completed_
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3401_request/$exit
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3401_request/ack
      -- 
    ack_7576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3401_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(465)); -- 
    -- CP-element group 466:  join  fork  transition  input  output  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	443 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	467 
    -- CP-element group 466:  members (24) 
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3401_update_completed_
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3401_complete/$exit
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3401_complete/ack
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_sample_start_
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_base_address_calculated
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_word_address_calculated
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_root_address_calculated
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_base_address_resized
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_base_addr_resize/$entry
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_base_addr_resize/$exit
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_base_addr_resize/base_resize_req
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_base_addr_resize/base_resize_ack
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_base_plus_offset/$entry
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_base_plus_offset/$exit
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_base_plus_offset/sum_rename_req
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_base_plus_offset/sum_rename_ack
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_word_addrgen/$entry
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_word_addrgen/$exit
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_word_addrgen/root_register_req
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_word_addrgen/root_register_ack
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Sample/$entry
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Sample/word_access_start/$entry
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Sample/word_access_start/word_0/$entry
      -- CP-element group 466: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Sample/word_access_start/word_0/rr
      -- 
    ack_7581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3401_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(466)); -- 
    rr_7614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(466), ack => ptr_deref_3405_load_0_req_0); -- 
    -- CP-element group 467:  transition  input  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	466 
    -- CP-element group 467: successors 
    -- CP-element group 467:  members (5) 
      -- CP-element group 467: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_sample_completed_
      -- CP-element group 467: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Sample/$exit
      -- CP-element group 467: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Sample/word_access_start/$exit
      -- CP-element group 467: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Sample/word_access_start/word_0/$exit
      -- CP-element group 467: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Sample/word_access_start/word_0/ra
      -- 
    ra_7615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3405_load_0_ack_0, ack => zeropad3D_CP_2152_elements(467)); -- 
    -- CP-element group 468:  transition  input  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	443 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	475 
    -- CP-element group 468:  members (9) 
      -- CP-element group 468: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_update_completed_
      -- CP-element group 468: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Update/$exit
      -- CP-element group 468: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Update/word_access_complete/$exit
      -- CP-element group 468: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Update/word_access_complete/word_0/$exit
      -- CP-element group 468: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Update/word_access_complete/word_0/ca
      -- CP-element group 468: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Update/ptr_deref_3405_Merge/$entry
      -- CP-element group 468: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Update/ptr_deref_3405_Merge/$exit
      -- CP-element group 468: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Update/ptr_deref_3405_Merge/merge_req
      -- CP-element group 468: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3405_Update/ptr_deref_3405_Merge/merge_ack
      -- 
    ca_7626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3405_load_0_ack_1, ack => zeropad3D_CP_2152_elements(468)); -- 
    -- CP-element group 469:  transition  input  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	460 
    -- CP-element group 469: successors 
    -- CP-element group 469:  members (3) 
      -- CP-element group 469: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3419_sample_completed_
      -- CP-element group 469: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3419_Sample/$exit
      -- CP-element group 469: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3419_Sample/ra
      -- 
    ra_7640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3419_inst_ack_0, ack => zeropad3D_CP_2152_elements(469)); -- 
    -- CP-element group 470:  transition  input  output  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	443 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	471 
    -- CP-element group 470:  members (16) 
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3419_update_completed_
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3419_Update/$exit
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/type_cast_3419_Update/ca
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_index_resized_1
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_index_scaled_1
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_index_computed_1
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_index_resize_1/$entry
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_index_resize_1/$exit
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_index_resize_1/index_resize_req
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_index_resize_1/index_resize_ack
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_index_scale_1/$entry
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_index_scale_1/$exit
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_index_scale_1/scale_rename_req
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_index_scale_1/scale_rename_ack
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_final_index_sum_regn_Sample/$entry
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_final_index_sum_regn_Sample/req
      -- 
    ca_7645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 470_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3419_inst_ack_1, ack => zeropad3D_CP_2152_elements(470)); -- 
    req_7670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(470), ack => array_obj_ref_3425_index_offset_req_0); -- 
    -- CP-element group 471:  transition  input  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	470 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	478 
    -- CP-element group 471:  members (3) 
      -- CP-element group 471: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_final_index_sum_regn_sample_complete
      -- CP-element group 471: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_final_index_sum_regn_Sample/$exit
      -- CP-element group 471: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_final_index_sum_regn_Sample/ack
      -- 
    ack_7671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3425_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(471)); -- 
    -- CP-element group 472:  transition  input  output  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	443 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	473 
    -- CP-element group 472:  members (11) 
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3426_request/req
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3426_request/$entry
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3426_sample_start_
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_root_address_calculated
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_offset_calculated
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_final_index_sum_regn_Update/$exit
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_final_index_sum_regn_Update/ack
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_base_plus_offset/$entry
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_base_plus_offset/$exit
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_base_plus_offset/sum_rename_req
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/array_obj_ref_3425_base_plus_offset/sum_rename_ack
      -- 
    ack_7676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3425_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(472)); -- 
    req_7685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(472), ack => addr_of_3426_final_reg_req_0); -- 
    -- CP-element group 473:  transition  input  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	472 
    -- CP-element group 473: successors 
    -- CP-element group 473:  members (3) 
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3426_request/ack
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3426_request/$exit
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3426_sample_completed_
      -- 
    ack_7686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3426_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(473)); -- 
    -- CP-element group 474:  fork  transition  input  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	443 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	475 
    -- CP-element group 474:  members (19) 
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_base_address_calculated
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_word_address_calculated
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_root_address_calculated
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_base_address_resized
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_base_addr_resize/$entry
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_base_addr_resize/$exit
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3426_complete/ack
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_word_addrgen/root_register_ack
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_word_addrgen/root_register_req
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_word_addrgen/$exit
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3426_complete/$exit
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_word_addrgen/$entry
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_base_plus_offset/sum_rename_ack
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_base_plus_offset/sum_rename_req
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_base_plus_offset/$exit
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_base_plus_offset/$entry
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_base_addr_resize/base_resize_ack
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_base_addr_resize/base_resize_req
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/addr_of_3426_update_completed_
      -- 
    ack_7691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 474_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3426_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(474)); -- 
    -- CP-element group 475:  join  transition  output  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	468 
    -- CP-element group 475: 	474 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	476 
    -- CP-element group 475:  members (9) 
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Sample/word_access_start/word_0/rr
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_sample_start_
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Sample/word_access_start/word_0/$entry
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Sample/word_access_start/$entry
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Sample/ptr_deref_3429_Split/split_ack
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Sample/ptr_deref_3429_Split/split_req
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Sample/ptr_deref_3429_Split/$exit
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Sample/ptr_deref_3429_Split/$entry
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Sample/$entry
      -- 
    rr_7729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(475), ack => ptr_deref_3429_store_0_req_0); -- 
    zeropad3D_cp_element_group_475: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_475"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(468) & zeropad3D_CP_2152_elements(474);
      gj_zeropad3D_cp_element_group_475 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(475), clk => clk, reset => reset); --
    end block;
    -- CP-element group 476:  transition  input  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	475 
    -- CP-element group 476: successors 
    -- CP-element group 476:  members (5) 
      -- CP-element group 476: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_sample_completed_
      -- CP-element group 476: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Sample/word_access_start/word_0/$exit
      -- CP-element group 476: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Sample/word_access_start/word_0/ra
      -- CP-element group 476: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Sample/word_access_start/$exit
      -- CP-element group 476: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Sample/$exit
      -- 
    ra_7730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 476_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3429_store_0_ack_0, ack => zeropad3D_CP_2152_elements(476)); -- 
    -- CP-element group 477:  transition  input  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	443 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	478 
    -- CP-element group 477:  members (5) 
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_update_completed_
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Update/$exit
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Update/word_access_complete/$exit
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Update/word_access_complete/word_0/ca
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/ptr_deref_3429_Update/word_access_complete/word_0/$exit
      -- 
    ca_7741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 477_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3429_store_0_ack_1, ack => zeropad3D_CP_2152_elements(477)); -- 
    -- CP-element group 478:  join  transition  place  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	463 
    -- CP-element group 478: 	471 
    -- CP-element group 478: 	477 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	1030 
    -- CP-element group 478:  members (5) 
      -- CP-element group 478: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431__exit__
      -- CP-element group 478: 	 branch_block_stmt_714/ifx_xelse956_ifx_xend1004
      -- CP-element group 478: 	 branch_block_stmt_714/assign_stmt_3331_to_assign_stmt_3431/$exit
      -- CP-element group 478: 	 branch_block_stmt_714/ifx_xelse956_ifx_xend1004_PhiReq/$entry
      -- CP-element group 478: 	 branch_block_stmt_714/ifx_xelse956_ifx_xend1004_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_478: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_478"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(463) & zeropad3D_CP_2152_elements(471) & zeropad3D_CP_2152_elements(477);
      gj_zeropad3D_cp_element_group_478 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(478), clk => clk, reset => reset); --
    end block;
    -- CP-element group 479:  transition  input  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	1030 
    -- CP-element group 479: successors 
    -- CP-element group 479:  members (3) 
      -- CP-element group 479: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/type_cast_3437_sample_completed_
      -- CP-element group 479: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/type_cast_3437_Sample/$exit
      -- CP-element group 479: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/type_cast_3437_Sample/ra
      -- 
    ra_7753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3437_inst_ack_0, ack => zeropad3D_CP_2152_elements(479)); -- 
    -- CP-element group 480:  branch  transition  place  input  output  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	1030 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	481 
    -- CP-element group 480: 	482 
    -- CP-element group 480:  members (13) 
      -- CP-element group 480: 	 branch_block_stmt_714/if_stmt_3452__entry__
      -- CP-element group 480: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451__exit__
      -- CP-element group 480: 	 branch_block_stmt_714/if_stmt_3452_eval_test/$entry
      -- CP-element group 480: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/type_cast_3437_update_completed_
      -- CP-element group 480: 	 branch_block_stmt_714/if_stmt_3452_eval_test/$exit
      -- CP-element group 480: 	 branch_block_stmt_714/if_stmt_3452_eval_test/branch_req
      -- CP-element group 480: 	 branch_block_stmt_714/if_stmt_3452_if_link/$entry
      -- CP-element group 480: 	 branch_block_stmt_714/if_stmt_3452_dead_link/$entry
      -- CP-element group 480: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/type_cast_3437_Update/ca
      -- CP-element group 480: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/$exit
      -- CP-element group 480: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/type_cast_3437_Update/$exit
      -- CP-element group 480: 	 branch_block_stmt_714/if_stmt_3452_else_link/$entry
      -- CP-element group 480: 	 branch_block_stmt_714/R_cmp1012_3453_place
      -- 
    ca_7758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 480_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3437_inst_ack_1, ack => zeropad3D_CP_2152_elements(480)); -- 
    branch_req_7766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(480), ack => if_stmt_3452_branch_req_0); -- 
    -- CP-element group 481:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	480 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	1039 
    -- CP-element group 481: 	1040 
    -- CP-element group 481: 	1042 
    -- CP-element group 481: 	1043 
    -- CP-element group 481: 	1045 
    -- CP-element group 481: 	1046 
    -- CP-element group 481:  members (40) 
      -- CP-element group 481: 	 branch_block_stmt_714/merge_stmt_3458__exit__
      -- CP-element group 481: 	 branch_block_stmt_714/assign_stmt_3464__entry__
      -- CP-element group 481: 	 branch_block_stmt_714/assign_stmt_3464__exit__
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057
      -- CP-element group 481: 	 branch_block_stmt_714/assign_stmt_3464/$exit
      -- CP-element group 481: 	 branch_block_stmt_714/assign_stmt_3464/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/if_stmt_3452_if_link/if_choice_transition
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xend1004_ifx_xthen1014
      -- CP-element group 481: 	 branch_block_stmt_714/if_stmt_3452_if_link/$exit
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xend1004_ifx_xthen1014_PhiReq/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xend1004_ifx_xthen1014_PhiReq/$exit
      -- CP-element group 481: 	 branch_block_stmt_714/merge_stmt_3458_PhiReqMerge
      -- CP-element group 481: 	 branch_block_stmt_714/merge_stmt_3458_PhiAck/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/merge_stmt_3458_PhiAck/$exit
      -- CP-element group 481: 	 branch_block_stmt_714/merge_stmt_3458_PhiAck/dummy
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/type_cast_3561/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/type_cast_3561/SplitProtocol/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/type_cast_3561/SplitProtocol/Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/type_cast_3561/SplitProtocol/Sample/rr
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/type_cast_3561/SplitProtocol/Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/type_cast_3561/SplitProtocol/Update/cr
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3568/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3568/SplitProtocol/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3568/SplitProtocol/Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3568/SplitProtocol/Sample/rr
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3568/SplitProtocol/Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3568/SplitProtocol/Update/cr
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3576/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3576/SplitProtocol/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3576/SplitProtocol/Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3576/SplitProtocol/Sample/rr
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3576/SplitProtocol/Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3576/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3452_branch_ack_1, ack => zeropad3D_CP_2152_elements(481)); -- 
    rr_12940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(481), ack => type_cast_3561_inst_req_0); -- 
    cr_12945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(481), ack => type_cast_3561_inst_req_1); -- 
    rr_12963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(481), ack => type_cast_3568_inst_req_0); -- 
    cr_12968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(481), ack => type_cast_3568_inst_req_1); -- 
    rr_12986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(481), ack => type_cast_3576_inst_req_0); -- 
    cr_12991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(481), ack => type_cast_3576_inst_req_1); -- 
    -- CP-element group 482:  fork  transition  place  input  output  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	480 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	483 
    -- CP-element group 482: 	484 
    -- CP-element group 482: 	485 
    -- CP-element group 482: 	486 
    -- CP-element group 482: 	488 
    -- CP-element group 482: 	491 
    -- CP-element group 482: 	493 
    -- CP-element group 482: 	494 
    -- CP-element group 482: 	495 
    -- CP-element group 482: 	497 
    -- CP-element group 482:  members (54) 
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550__entry__
      -- CP-element group 482: 	 branch_block_stmt_714/merge_stmt_3466__exit__
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3503_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Update/word_access_complete/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Update/word_access_complete/word_0/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3527_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Update/word_access_complete/word_0/cr
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3520_update_start_
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Update/word_access_complete/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3527_update_start_
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Update/word_access_complete/word_0/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Sample/word_access_start/word_0/rr
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Sample/word_access_start/word_0/rr
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3503_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Sample/word_access_start/word_0/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Sample/word_access_start/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Sample/word_access_start/word_0/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3503_update_start_
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3483_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_root_address_calculated
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Sample/word_access_start/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3527_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_root_address_calculated
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_word_address_calculated
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_update_start_
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3476_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_word_address_calculated
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_update_start_
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3476_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3483_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3476_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3520_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3520_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3476_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3476_update_start_
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3476_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/ifx_xend1004_ifx_xelse1019
      -- CP-element group 482: 	 branch_block_stmt_714/if_stmt_3452_else_link/else_choice_transition
      -- CP-element group 482: 	 branch_block_stmt_714/if_stmt_3452_else_link/$exit
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Update/word_access_complete/word_0/cr
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3483_update_start_
      -- CP-element group 482: 	 branch_block_stmt_714/ifx_xend1004_ifx_xelse1019_PhiReq/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/ifx_xend1004_ifx_xelse1019_PhiReq/$exit
      -- CP-element group 482: 	 branch_block_stmt_714/merge_stmt_3466_PhiReqMerge
      -- CP-element group 482: 	 branch_block_stmt_714/merge_stmt_3466_PhiAck/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/merge_stmt_3466_PhiAck/$exit
      -- CP-element group 482: 	 branch_block_stmt_714/merge_stmt_3466_PhiAck/dummy
      -- 
    else_choice_transition_7775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 482_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3452_branch_ack_0, ack => zeropad3D_CP_2152_elements(482)); -- 
    cr_7857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(482), ack => type_cast_3503_inst_req_1); -- 
    cr_7918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(482), ack => type_cast_3527_inst_req_1); -- 
    cr_7824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(482), ack => LOAD_col_high_3479_load_0_req_1); -- 
    rr_7813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(482), ack => LOAD_col_high_3479_load_0_req_0); -- 
    rr_7888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(482), ack => LOAD_row_high_3523_load_0_req_0); -- 
    cr_7843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(482), ack => type_cast_3483_inst_req_1); -- 
    cr_7796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(482), ack => type_cast_3476_inst_req_1); -- 
    rr_7791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(482), ack => type_cast_3476_inst_req_0); -- 
    cr_7871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(482), ack => type_cast_3520_inst_req_1); -- 
    cr_7899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(482), ack => LOAD_row_high_3523_load_0_req_1); -- 
    -- CP-element group 483:  transition  input  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	482 
    -- CP-element group 483: successors 
    -- CP-element group 483:  members (3) 
      -- CP-element group 483: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3476_Sample/ra
      -- CP-element group 483: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3476_Sample/$exit
      -- CP-element group 483: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3476_sample_completed_
      -- 
    ra_7792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 483_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3476_inst_ack_0, ack => zeropad3D_CP_2152_elements(483)); -- 
    -- CP-element group 484:  transition  input  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	482 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	489 
    -- CP-element group 484:  members (3) 
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3476_Update/ca
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3476_Update/$exit
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3476_update_completed_
      -- 
    ca_7797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3476_inst_ack_1, ack => zeropad3D_CP_2152_elements(484)); -- 
    -- CP-element group 485:  transition  input  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	482 
    -- CP-element group 485: successors 
    -- CP-element group 485:  members (5) 
      -- CP-element group 485: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Sample/word_access_start/word_0/ra
      -- CP-element group 485: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Sample/word_access_start/word_0/$exit
      -- CP-element group 485: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Sample/word_access_start/$exit
      -- CP-element group 485: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Sample/$exit
      -- CP-element group 485: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_sample_completed_
      -- 
    ra_7814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3479_load_0_ack_0, ack => zeropad3D_CP_2152_elements(485)); -- 
    -- CP-element group 486:  transition  input  output  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	482 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	487 
    -- CP-element group 486:  members (12) 
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Update/$exit
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Update/word_access_complete/$exit
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Update/word_access_complete/word_0/$exit
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Update/word_access_complete/word_0/ca
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Update/LOAD_col_high_3479_Merge/$entry
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Update/LOAD_col_high_3479_Merge/$exit
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Update/LOAD_col_high_3479_Merge/merge_req
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_Update/LOAD_col_high_3479_Merge/merge_ack
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_col_high_3479_update_completed_
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3483_Sample/rr
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3483_Sample/$entry
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3483_sample_start_
      -- 
    ca_7825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 486_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3479_load_0_ack_1, ack => zeropad3D_CP_2152_elements(486)); -- 
    rr_7838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(486), ack => type_cast_3483_inst_req_0); -- 
    -- CP-element group 487:  transition  input  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	486 
    -- CP-element group 487: successors 
    -- CP-element group 487:  members (3) 
      -- CP-element group 487: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3483_Sample/ra
      -- CP-element group 487: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3483_Sample/$exit
      -- CP-element group 487: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3483_sample_completed_
      -- 
    ra_7839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 487_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3483_inst_ack_0, ack => zeropad3D_CP_2152_elements(487)); -- 
    -- CP-element group 488:  transition  input  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	482 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	489 
    -- CP-element group 488:  members (3) 
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3483_Update/ca
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3483_Update/$exit
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3483_update_completed_
      -- 
    ca_7844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3483_inst_ack_1, ack => zeropad3D_CP_2152_elements(488)); -- 
    -- CP-element group 489:  join  transition  output  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	484 
    -- CP-element group 489: 	488 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	490 
    -- CP-element group 489:  members (3) 
      -- CP-element group 489: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3503_Sample/rr
      -- CP-element group 489: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3503_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3503_sample_start_
      -- 
    rr_7852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(489), ack => type_cast_3503_inst_req_0); -- 
    zeropad3D_cp_element_group_489: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_489"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(484) & zeropad3D_CP_2152_elements(488);
      gj_zeropad3D_cp_element_group_489 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(489), clk => clk, reset => reset); --
    end block;
    -- CP-element group 490:  transition  input  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	489 
    -- CP-element group 490: successors 
    -- CP-element group 490:  members (3) 
      -- CP-element group 490: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3503_Sample/$exit
      -- CP-element group 490: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3503_Sample/ra
      -- CP-element group 490: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3503_sample_completed_
      -- 
    ra_7853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 490_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3503_inst_ack_0, ack => zeropad3D_CP_2152_elements(490)); -- 
    -- CP-element group 491:  transition  input  output  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	482 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	492 
    -- CP-element group 491:  members (6) 
      -- CP-element group 491: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3503_Update/$exit
      -- CP-element group 491: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3503_Update/ca
      -- CP-element group 491: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3520_sample_start_
      -- CP-element group 491: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3503_update_completed_
      -- CP-element group 491: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3520_Sample/rr
      -- CP-element group 491: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3520_Sample/$entry
      -- 
    ca_7858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3503_inst_ack_1, ack => zeropad3D_CP_2152_elements(491)); -- 
    rr_7866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(491), ack => type_cast_3520_inst_req_0); -- 
    -- CP-element group 492:  transition  input  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	491 
    -- CP-element group 492: successors 
    -- CP-element group 492:  members (3) 
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3520_sample_completed_
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3520_Sample/ra
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3520_Sample/$exit
      -- 
    ra_7867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3520_inst_ack_0, ack => zeropad3D_CP_2152_elements(492)); -- 
    -- CP-element group 493:  transition  input  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	482 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	498 
    -- CP-element group 493:  members (3) 
      -- CP-element group 493: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3520_Update/ca
      -- CP-element group 493: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3520_Update/$exit
      -- CP-element group 493: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3520_update_completed_
      -- 
    ca_7872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 493_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3520_inst_ack_1, ack => zeropad3D_CP_2152_elements(493)); -- 
    -- CP-element group 494:  transition  input  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	482 
    -- CP-element group 494: successors 
    -- CP-element group 494:  members (5) 
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Sample/word_access_start/word_0/ra
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Sample/word_access_start/word_0/$exit
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Sample/word_access_start/$exit
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Sample/$exit
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_sample_completed_
      -- 
    ra_7889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 494_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3523_load_0_ack_0, ack => zeropad3D_CP_2152_elements(494)); -- 
    -- CP-element group 495:  transition  input  output  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	482 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	496 
    -- CP-element group 495:  members (12) 
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Update/LOAD_row_high_3523_Merge/merge_ack
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Update/$exit
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3527_Sample/$entry
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3527_sample_start_
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Update/word_access_complete/$exit
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Update/word_access_complete/word_0/$exit
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Update/LOAD_row_high_3523_Merge/merge_req
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Update/LOAD_row_high_3523_Merge/$exit
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Update/LOAD_row_high_3523_Merge/$entry
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_update_completed_
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/LOAD_row_high_3523_Update/word_access_complete/word_0/ca
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3527_Sample/rr
      -- 
    ca_7900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3523_load_0_ack_1, ack => zeropad3D_CP_2152_elements(495)); -- 
    rr_7913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(495), ack => type_cast_3527_inst_req_0); -- 
    -- CP-element group 496:  transition  input  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	495 
    -- CP-element group 496: successors 
    -- CP-element group 496:  members (3) 
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3527_Sample/$exit
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3527_sample_completed_
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3527_Sample/ra
      -- 
    ra_7914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 496_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3527_inst_ack_0, ack => zeropad3D_CP_2152_elements(496)); -- 
    -- CP-element group 497:  transition  input  bypass 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	482 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	498 
    -- CP-element group 497:  members (3) 
      -- CP-element group 497: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3527_Update/ca
      -- CP-element group 497: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3527_Update/$exit
      -- CP-element group 497: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/type_cast_3527_update_completed_
      -- 
    ca_7919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 497_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3527_inst_ack_1, ack => zeropad3D_CP_2152_elements(497)); -- 
    -- CP-element group 498:  branch  join  transition  place  output  bypass 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	493 
    -- CP-element group 498: 	497 
    -- CP-element group 498: successors 
    -- CP-element group 498: 	499 
    -- CP-element group 498: 	500 
    -- CP-element group 498:  members (10) 
      -- CP-element group 498: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550__exit__
      -- CP-element group 498: 	 branch_block_stmt_714/if_stmt_3551__entry__
      -- CP-element group 498: 	 branch_block_stmt_714/if_stmt_3551_dead_link/$entry
      -- CP-element group 498: 	 branch_block_stmt_714/if_stmt_3551_else_link/$entry
      -- CP-element group 498: 	 branch_block_stmt_714/R_cmp1048_3552_place
      -- CP-element group 498: 	 branch_block_stmt_714/assign_stmt_3472_to_assign_stmt_3550/$exit
      -- CP-element group 498: 	 branch_block_stmt_714/if_stmt_3551_if_link/$entry
      -- CP-element group 498: 	 branch_block_stmt_714/if_stmt_3551_eval_test/branch_req
      -- CP-element group 498: 	 branch_block_stmt_714/if_stmt_3551_eval_test/$exit
      -- CP-element group 498: 	 branch_block_stmt_714/if_stmt_3551_eval_test/$entry
      -- 
    branch_req_7927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(498), ack => if_stmt_3551_branch_req_0); -- 
    zeropad3D_cp_element_group_498: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_498"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(493) & zeropad3D_CP_2152_elements(497);
      gj_zeropad3D_cp_element_group_498 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(498), clk => clk, reset => reset); --
    end block;
    -- CP-element group 499:  fork  transition  place  input  output  bypass 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	498 
    -- CP-element group 499: successors 
    -- CP-element group 499: 	1054 
    -- CP-element group 499: 	1055 
    -- CP-element group 499: 	1057 
    -- CP-element group 499: 	1058 
    -- CP-element group 499: 	1060 
    -- CP-element group 499: 	1061 
    -- CP-element group 499:  members (28) 
      -- CP-element group 499: 	 branch_block_stmt_714/if_stmt_3551_if_link/if_choice_transition
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058
      -- CP-element group 499: 	 branch_block_stmt_714/if_stmt_3551_if_link/$exit
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/type_cast_3583/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/type_cast_3583/SplitProtocol/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/type_cast_3583/SplitProtocol/Sample/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/type_cast_3583/SplitProtocol/Sample/rr
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/type_cast_3583/SplitProtocol/Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/type_cast_3583/SplitProtocol/Update/cr
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/type_cast_3587/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/type_cast_3587/SplitProtocol/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/type_cast_3587/SplitProtocol/Sample/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/type_cast_3587/SplitProtocol/Sample/rr
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/type_cast_3587/SplitProtocol/Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/type_cast_3587/SplitProtocol/Update/cr
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/type_cast_3591/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/type_cast_3591/SplitProtocol/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/type_cast_3591/SplitProtocol/Sample/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/type_cast_3591/SplitProtocol/Sample/rr
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/type_cast_3591/SplitProtocol/Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/type_cast_3591/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 499_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3551_branch_ack_1, ack => zeropad3D_CP_2152_elements(499)); -- 
    rr_13019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(499), ack => type_cast_3583_inst_req_0); -- 
    cr_13024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(499), ack => type_cast_3583_inst_req_1); -- 
    rr_13042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(499), ack => type_cast_3587_inst_req_0); -- 
    cr_13047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(499), ack => type_cast_3587_inst_req_1); -- 
    rr_13065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(499), ack => type_cast_3591_inst_req_0); -- 
    cr_13070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(499), ack => type_cast_3591_inst_req_1); -- 
    -- CP-element group 500:  fork  transition  place  input  output  bypass 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	498 
    -- CP-element group 500: successors 
    -- CP-element group 500: 	1031 
    -- CP-element group 500: 	1032 
    -- CP-element group 500: 	1033 
    -- CP-element group 500: 	1035 
    -- CP-element group 500: 	1036 
    -- CP-element group 500:  members (22) 
      -- CP-element group 500: 	 branch_block_stmt_714/if_stmt_3551_else_link/else_choice_transition
      -- CP-element group 500: 	 branch_block_stmt_714/if_stmt_3551_else_link/$exit
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3558/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3570/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3570/SplitProtocol/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3570/SplitProtocol/Sample/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3570/SplitProtocol/Sample/rr
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3570/SplitProtocol/Update/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3570/SplitProtocol/Update/cr
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3574/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3574/SplitProtocol/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3574/SplitProtocol/Sample/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3574/SplitProtocol/Sample/rr
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3574/SplitProtocol/Update/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3574/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 500_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3551_branch_ack_0, ack => zeropad3D_CP_2152_elements(500)); -- 
    rr_12891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(500), ack => type_cast_3570_inst_req_0); -- 
    cr_12896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(500), ack => type_cast_3570_inst_req_1); -- 
    rr_12914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(500), ack => type_cast_3574_inst_req_0); -- 
    cr_12919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(500), ack => type_cast_3574_inst_req_1); -- 
    -- CP-element group 501:  transition  input  bypass 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	1067 
    -- CP-element group 501: successors 
    -- CP-element group 501:  members (3) 
      -- CP-element group 501: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3595_Sample/$exit
      -- CP-element group 501: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3595_Sample/ra
      -- CP-element group 501: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3595_sample_completed_
      -- 
    ra_7950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 501_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3595_inst_ack_0, ack => zeropad3D_CP_2152_elements(501)); -- 
    -- CP-element group 502:  transition  input  bypass 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	1067 
    -- CP-element group 502: successors 
    -- CP-element group 502: 	517 
    -- CP-element group 502:  members (3) 
      -- CP-element group 502: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3595_Update/$exit
      -- CP-element group 502: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3595_Update/ca
      -- CP-element group 502: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3595_update_completed_
      -- 
    ca_7955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 502_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3595_inst_ack_1, ack => zeropad3D_CP_2152_elements(502)); -- 
    -- CP-element group 503:  transition  input  bypass 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	1067 
    -- CP-element group 503: successors 
    -- CP-element group 503:  members (3) 
      -- CP-element group 503: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3605_Sample/ra
      -- CP-element group 503: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3605_Sample/$exit
      -- CP-element group 503: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3605_sample_completed_
      -- 
    ra_7964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 503_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3605_inst_ack_0, ack => zeropad3D_CP_2152_elements(503)); -- 
    -- CP-element group 504:  transition  input  bypass 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: 	1067 
    -- CP-element group 504: successors 
    -- CP-element group 504: 	517 
    -- CP-element group 504:  members (3) 
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3605_Update/$exit
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3605_Update/ca
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3605_update_completed_
      -- 
    ca_7969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 504_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3605_inst_ack_1, ack => zeropad3D_CP_2152_elements(504)); -- 
    -- CP-element group 505:  transition  input  bypass 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	1067 
    -- CP-element group 505: successors 
    -- CP-element group 505:  members (5) 
      -- CP-element group 505: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_sample_completed_
      -- CP-element group 505: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Sample/$exit
      -- CP-element group 505: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Sample/word_access_start/$exit
      -- CP-element group 505: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Sample/word_access_start/word_0/$exit
      -- CP-element group 505: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Sample/word_access_start/word_0/ra
      -- 
    ra_7986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 505_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3614_load_0_ack_0, ack => zeropad3D_CP_2152_elements(505)); -- 
    -- CP-element group 506:  transition  input  output  bypass 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	1067 
    -- CP-element group 506: successors 
    -- CP-element group 506: 	515 
    -- CP-element group 506:  members (12) 
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_update_completed_
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Update/$exit
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Update/word_access_complete/$exit
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Update/word_access_complete/word_0/$exit
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Update/word_access_complete/word_0/ca
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Update/LOAD_pad_3614_Merge/$entry
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Update/LOAD_pad_3614_Merge/$exit
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Update/LOAD_pad_3614_Merge/merge_req
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Update/LOAD_pad_3614_Merge/merge_ack
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3684_sample_start_
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3684_Sample/$entry
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3684_Sample/rr
      -- 
    ca_7997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 506_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3614_load_0_ack_1, ack => zeropad3D_CP_2152_elements(506)); -- 
    rr_8157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(506), ack => type_cast_3684_inst_req_0); -- 
    -- CP-element group 507:  transition  input  bypass 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	1067 
    -- CP-element group 507: successors 
    -- CP-element group 507:  members (5) 
      -- CP-element group 507: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_sample_completed_
      -- CP-element group 507: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Sample/$exit
      -- CP-element group 507: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Sample/word_access_start/$exit
      -- CP-element group 507: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Sample/word_access_start/word_0/$exit
      -- CP-element group 507: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Sample/word_access_start/word_0/ra
      -- 
    ra_8019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 507_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_3617_load_0_ack_0, ack => zeropad3D_CP_2152_elements(507)); -- 
    -- CP-element group 508:  transition  input  output  bypass 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: 	1067 
    -- CP-element group 508: successors 
    -- CP-element group 508: 	513 
    -- CP-element group 508:  members (12) 
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_update_completed_
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Update/$exit
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Update/word_access_complete/$exit
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Update/word_access_complete/word_0/$exit
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Update/word_access_complete/word_0/ca
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Update/LOAD_depth_high_3617_Merge/$entry
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Update/LOAD_depth_high_3617_Merge/$exit
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Update/LOAD_depth_high_3617_Merge/merge_req
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Update/LOAD_depth_high_3617_Merge/merge_ack
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3645_sample_start_
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3645_Sample/$entry
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3645_Sample/rr
      -- 
    ca_8030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 508_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_3617_load_0_ack_1, ack => zeropad3D_CP_2152_elements(508)); -- 
    rr_8143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(508), ack => type_cast_3645_inst_req_0); -- 
    -- CP-element group 509:  transition  input  bypass 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	1067 
    -- CP-element group 509: successors 
    -- CP-element group 509:  members (5) 
      -- CP-element group 509: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_sample_completed_
      -- CP-element group 509: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Sample/$exit
      -- CP-element group 509: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Sample/word_access_start/$exit
      -- CP-element group 509: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Sample/word_access_start/word_0/$exit
      -- CP-element group 509: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Sample/word_access_start/word_0/ra
      -- 
    ra_8069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 509_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3629_load_0_ack_0, ack => zeropad3D_CP_2152_elements(509)); -- 
    -- CP-element group 510:  transition  input  bypass 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	1067 
    -- CP-element group 510: successors 
    -- CP-element group 510: 	517 
    -- CP-element group 510:  members (9) 
      -- CP-element group 510: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_update_completed_
      -- CP-element group 510: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Update/$exit
      -- CP-element group 510: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Update/word_access_complete/$exit
      -- CP-element group 510: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Update/word_access_complete/word_0/$exit
      -- CP-element group 510: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Update/word_access_complete/word_0/ca
      -- CP-element group 510: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Update/ptr_deref_3629_Merge/$entry
      -- CP-element group 510: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Update/ptr_deref_3629_Merge/$exit
      -- CP-element group 510: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Update/ptr_deref_3629_Merge/merge_req
      -- CP-element group 510: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Update/ptr_deref_3629_Merge/merge_ack
      -- 
    ca_8080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 510_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3629_load_0_ack_1, ack => zeropad3D_CP_2152_elements(510)); -- 
    -- CP-element group 511:  transition  input  bypass 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	1067 
    -- CP-element group 511: successors 
    -- CP-element group 511:  members (5) 
      -- CP-element group 511: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_sample_completed_
      -- CP-element group 511: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Sample/$exit
      -- CP-element group 511: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Sample/word_access_start/$exit
      -- CP-element group 511: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Sample/word_access_start/word_0/$exit
      -- CP-element group 511: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Sample/word_access_start/word_0/ra
      -- 
    ra_8119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 511_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3641_load_0_ack_0, ack => zeropad3D_CP_2152_elements(511)); -- 
    -- CP-element group 512:  transition  input  bypass 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: 	1067 
    -- CP-element group 512: successors 
    -- CP-element group 512: 	517 
    -- CP-element group 512:  members (9) 
      -- CP-element group 512: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_update_completed_
      -- CP-element group 512: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Update/$exit
      -- CP-element group 512: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Update/word_access_complete/$exit
      -- CP-element group 512: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Update/word_access_complete/word_0/$exit
      -- CP-element group 512: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Update/word_access_complete/word_0/ca
      -- CP-element group 512: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Update/ptr_deref_3641_Merge/$entry
      -- CP-element group 512: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Update/ptr_deref_3641_Merge/$exit
      -- CP-element group 512: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Update/ptr_deref_3641_Merge/merge_req
      -- CP-element group 512: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Update/ptr_deref_3641_Merge/merge_ack
      -- 
    ca_8130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 512_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3641_load_0_ack_1, ack => zeropad3D_CP_2152_elements(512)); -- 
    -- CP-element group 513:  transition  input  bypass 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	508 
    -- CP-element group 513: successors 
    -- CP-element group 513:  members (3) 
      -- CP-element group 513: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3645_sample_completed_
      -- CP-element group 513: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3645_Sample/$exit
      -- CP-element group 513: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3645_Sample/ra
      -- 
    ra_8144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 513_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3645_inst_ack_0, ack => zeropad3D_CP_2152_elements(513)); -- 
    -- CP-element group 514:  transition  input  bypass 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	1067 
    -- CP-element group 514: successors 
    -- CP-element group 514: 	517 
    -- CP-element group 514:  members (3) 
      -- CP-element group 514: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3645_update_completed_
      -- CP-element group 514: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3645_Update/$exit
      -- CP-element group 514: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3645_Update/ca
      -- 
    ca_8149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 514_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3645_inst_ack_1, ack => zeropad3D_CP_2152_elements(514)); -- 
    -- CP-element group 515:  transition  input  bypass 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	506 
    -- CP-element group 515: successors 
    -- CP-element group 515:  members (3) 
      -- CP-element group 515: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3684_sample_completed_
      -- CP-element group 515: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3684_Sample/$exit
      -- CP-element group 515: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3684_Sample/ra
      -- 
    ra_8158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 515_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3684_inst_ack_0, ack => zeropad3D_CP_2152_elements(515)); -- 
    -- CP-element group 516:  transition  input  bypass 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: 	1067 
    -- CP-element group 516: successors 
    -- CP-element group 516: 	517 
    -- CP-element group 516:  members (3) 
      -- CP-element group 516: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3684_update_completed_
      -- CP-element group 516: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3684_Update/$exit
      -- CP-element group 516: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3684_Update/ca
      -- 
    ca_8163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 516_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3684_inst_ack_1, ack => zeropad3D_CP_2152_elements(516)); -- 
    -- CP-element group 517:  join  fork  transition  place  output  bypass 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	502 
    -- CP-element group 517: 	504 
    -- CP-element group 517: 	510 
    -- CP-element group 517: 	512 
    -- CP-element group 517: 	514 
    -- CP-element group 517: 	516 
    -- CP-element group 517: successors 
    -- CP-element group 517: 	1078 
    -- CP-element group 517: 	1079 
    -- CP-element group 517: 	1080 
    -- CP-element group 517: 	1082 
    -- CP-element group 517: 	1083 
    -- CP-element group 517:  members (22) 
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726__exit__
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/$exit
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3729/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3741/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3741/SplitProtocol/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3741/SplitProtocol/Sample/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3741/SplitProtocol/Sample/rr
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3741/SplitProtocol/Update/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3741/SplitProtocol/Update/cr
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3745/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3745/SplitProtocol/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3745/SplitProtocol/Sample/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3745/SplitProtocol/Sample/rr
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3745/SplitProtocol/Update/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3745/SplitProtocol/Update/cr
      -- 
    rr_13178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(517), ack => type_cast_3741_inst_req_0); -- 
    cr_13183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(517), ack => type_cast_3741_inst_req_1); -- 
    rr_13201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(517), ack => type_cast_3745_inst_req_0); -- 
    cr_13206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(517), ack => type_cast_3745_inst_req_1); -- 
    zeropad3D_cp_element_group_517: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_517"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(502) & zeropad3D_CP_2152_elements(504) & zeropad3D_CP_2152_elements(510) & zeropad3D_CP_2152_elements(512) & zeropad3D_CP_2152_elements(514) & zeropad3D_CP_2152_elements(516);
      gj_zeropad3D_cp_element_group_517 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(517), clk => clk, reset => reset); --
    end block;
    -- CP-element group 518:  transition  input  bypass 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	1090 
    -- CP-element group 518: successors 
    -- CP-element group 518:  members (3) 
      -- CP-element group 518: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/type_cast_3752_sample_completed_
      -- CP-element group 518: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/type_cast_3752_Sample/$exit
      -- CP-element group 518: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/type_cast_3752_Sample/ra
      -- 
    ra_8175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 518_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3752_inst_ack_0, ack => zeropad3D_CP_2152_elements(518)); -- 
    -- CP-element group 519:  branch  transition  place  input  output  bypass 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	1090 
    -- CP-element group 519: successors 
    -- CP-element group 519: 	520 
    -- CP-element group 519: 	521 
    -- CP-element group 519:  members (13) 
      -- CP-element group 519: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760__exit__
      -- CP-element group 519: 	 branch_block_stmt_714/if_stmt_3761__entry__
      -- CP-element group 519: 	 branch_block_stmt_714/R_cmp1127_3762_place
      -- CP-element group 519: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/$exit
      -- CP-element group 519: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/type_cast_3752_update_completed_
      -- CP-element group 519: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/type_cast_3752_Update/$exit
      -- CP-element group 519: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/type_cast_3752_Update/ca
      -- CP-element group 519: 	 branch_block_stmt_714/if_stmt_3761_dead_link/$entry
      -- CP-element group 519: 	 branch_block_stmt_714/if_stmt_3761_eval_test/$entry
      -- CP-element group 519: 	 branch_block_stmt_714/if_stmt_3761_eval_test/$exit
      -- CP-element group 519: 	 branch_block_stmt_714/if_stmt_3761_eval_test/branch_req
      -- CP-element group 519: 	 branch_block_stmt_714/if_stmt_3761_if_link/$entry
      -- CP-element group 519: 	 branch_block_stmt_714/if_stmt_3761_else_link/$entry
      -- 
    ca_8180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 519_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3752_inst_ack_1, ack => zeropad3D_CP_2152_elements(519)); -- 
    branch_req_8188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(519), ack => if_stmt_3761_branch_req_0); -- 
    -- CP-element group 520:  transition  place  input  bypass 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: 	519 
    -- CP-element group 520: successors 
    -- CP-element group 520: 	1091 
    -- CP-element group 520:  members (5) 
      -- CP-element group 520: 	 branch_block_stmt_714/whilex_xbody1122_ifx_xthen1158
      -- CP-element group 520: 	 branch_block_stmt_714/if_stmt_3761_if_link/$exit
      -- CP-element group 520: 	 branch_block_stmt_714/if_stmt_3761_if_link/if_choice_transition
      -- CP-element group 520: 	 branch_block_stmt_714/whilex_xbody1122_ifx_xthen1158_PhiReq/$entry
      -- CP-element group 520: 	 branch_block_stmt_714/whilex_xbody1122_ifx_xthen1158_PhiReq/$exit
      -- 
    if_choice_transition_8193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 520_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3761_branch_ack_1, ack => zeropad3D_CP_2152_elements(520)); -- 
    -- CP-element group 521:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	519 
    -- CP-element group 521: successors 
    -- CP-element group 521: 	522 
    -- CP-element group 521: 	523 
    -- CP-element group 521: 	525 
    -- CP-element group 521:  members (27) 
      -- CP-element group 521: 	 branch_block_stmt_714/merge_stmt_3767__exit__
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798__entry__
      -- CP-element group 521: 	 branch_block_stmt_714/whilex_xbody1122_lorx_xlhsx_xfalse1129
      -- CP-element group 521: 	 branch_block_stmt_714/if_stmt_3761_else_link/$exit
      -- CP-element group 521: 	 branch_block_stmt_714/if_stmt_3761_else_link/else_choice_transition
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_sample_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_update_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_word_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_root_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Sample/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Sample/word_access_start/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Sample/word_access_start/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Sample/word_access_start/word_0/rr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Update/word_access_complete/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Update/word_access_complete/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Update/word_access_complete/word_0/cr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/type_cast_3773_update_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/type_cast_3773_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/type_cast_3773_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_714/whilex_xbody1122_lorx_xlhsx_xfalse1129_PhiReq/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/whilex_xbody1122_lorx_xlhsx_xfalse1129_PhiReq/$exit
      -- CP-element group 521: 	 branch_block_stmt_714/merge_stmt_3767_PhiReqMerge
      -- CP-element group 521: 	 branch_block_stmt_714/merge_stmt_3767_PhiAck/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/merge_stmt_3767_PhiAck/$exit
      -- CP-element group 521: 	 branch_block_stmt_714/merge_stmt_3767_PhiAck/dummy
      -- 
    else_choice_transition_8197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 521_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3761_branch_ack_0, ack => zeropad3D_CP_2152_elements(521)); -- 
    rr_8218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => LOAD_row_high_3769_load_0_req_0); -- 
    cr_8229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => LOAD_row_high_3769_load_0_req_1); -- 
    cr_8248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => type_cast_3773_inst_req_1); -- 
    -- CP-element group 522:  transition  input  bypass 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	521 
    -- CP-element group 522: successors 
    -- CP-element group 522:  members (5) 
      -- CP-element group 522: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_sample_completed_
      -- CP-element group 522: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Sample/$exit
      -- CP-element group 522: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Sample/word_access_start/$exit
      -- CP-element group 522: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Sample/word_access_start/word_0/$exit
      -- CP-element group 522: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Sample/word_access_start/word_0/ra
      -- 
    ra_8219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 522_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3769_load_0_ack_0, ack => zeropad3D_CP_2152_elements(522)); -- 
    -- CP-element group 523:  transition  input  output  bypass 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: 	521 
    -- CP-element group 523: successors 
    -- CP-element group 523: 	524 
    -- CP-element group 523:  members (12) 
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_update_completed_
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Update/$exit
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Update/word_access_complete/$exit
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Update/word_access_complete/word_0/$exit
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Update/word_access_complete/word_0/ca
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Update/LOAD_row_high_3769_Merge/$entry
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Update/LOAD_row_high_3769_Merge/$exit
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Update/LOAD_row_high_3769_Merge/merge_req
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/LOAD_row_high_3769_Update/LOAD_row_high_3769_Merge/merge_ack
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/type_cast_3773_sample_start_
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/type_cast_3773_Sample/$entry
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/type_cast_3773_Sample/rr
      -- 
    ca_8230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 523_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3769_load_0_ack_1, ack => zeropad3D_CP_2152_elements(523)); -- 
    rr_8243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(523), ack => type_cast_3773_inst_req_0); -- 
    -- CP-element group 524:  transition  input  bypass 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: 	523 
    -- CP-element group 524: successors 
    -- CP-element group 524:  members (3) 
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/type_cast_3773_sample_completed_
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/type_cast_3773_Sample/$exit
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/type_cast_3773_Sample/ra
      -- 
    ra_8244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 524_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3773_inst_ack_0, ack => zeropad3D_CP_2152_elements(524)); -- 
    -- CP-element group 525:  branch  transition  place  input  output  bypass 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	521 
    -- CP-element group 525: successors 
    -- CP-element group 525: 	526 
    -- CP-element group 525: 	527 
    -- CP-element group 525:  members (13) 
      -- CP-element group 525: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798__exit__
      -- CP-element group 525: 	 branch_block_stmt_714/if_stmt_3799__entry__
      -- CP-element group 525: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/$exit
      -- CP-element group 525: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/type_cast_3773_update_completed_
      -- CP-element group 525: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/type_cast_3773_Update/$exit
      -- CP-element group 525: 	 branch_block_stmt_714/assign_stmt_3770_to_assign_stmt_3798/type_cast_3773_Update/ca
      -- CP-element group 525: 	 branch_block_stmt_714/if_stmt_3799_dead_link/$entry
      -- CP-element group 525: 	 branch_block_stmt_714/if_stmt_3799_eval_test/$entry
      -- CP-element group 525: 	 branch_block_stmt_714/if_stmt_3799_eval_test/$exit
      -- CP-element group 525: 	 branch_block_stmt_714/if_stmt_3799_eval_test/branch_req
      -- CP-element group 525: 	 branch_block_stmt_714/R_cmp1139_3800_place
      -- CP-element group 525: 	 branch_block_stmt_714/if_stmt_3799_if_link/$entry
      -- CP-element group 525: 	 branch_block_stmt_714/if_stmt_3799_else_link/$entry
      -- 
    ca_8249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 525_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3773_inst_ack_1, ack => zeropad3D_CP_2152_elements(525)); -- 
    branch_req_8257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(525), ack => if_stmt_3799_branch_req_0); -- 
    -- CP-element group 526:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: 	525 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	528 
    -- CP-element group 526: 	529 
    -- CP-element group 526:  members (18) 
      -- CP-element group 526: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817__entry__
      -- CP-element group 526: 	 branch_block_stmt_714/merge_stmt_3805__exit__
      -- CP-element group 526: 	 branch_block_stmt_714/if_stmt_3799_if_link/$exit
      -- CP-element group 526: 	 branch_block_stmt_714/if_stmt_3799_if_link/if_choice_transition
      -- CP-element group 526: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1129_lorx_xlhsx_xfalse1141
      -- CP-element group 526: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/$entry
      -- CP-element group 526: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/type_cast_3809_sample_start_
      -- CP-element group 526: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/type_cast_3809_update_start_
      -- CP-element group 526: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/type_cast_3809_Sample/$entry
      -- CP-element group 526: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/type_cast_3809_Sample/rr
      -- CP-element group 526: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/type_cast_3809_Update/$entry
      -- CP-element group 526: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/type_cast_3809_Update/cr
      -- CP-element group 526: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1129_lorx_xlhsx_xfalse1141_PhiReq/$entry
      -- CP-element group 526: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1129_lorx_xlhsx_xfalse1141_PhiReq/$exit
      -- CP-element group 526: 	 branch_block_stmt_714/merge_stmt_3805_PhiReqMerge
      -- CP-element group 526: 	 branch_block_stmt_714/merge_stmt_3805_PhiAck/$entry
      -- CP-element group 526: 	 branch_block_stmt_714/merge_stmt_3805_PhiAck/$exit
      -- CP-element group 526: 	 branch_block_stmt_714/merge_stmt_3805_PhiAck/dummy
      -- 
    if_choice_transition_8262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 526_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3799_branch_ack_1, ack => zeropad3D_CP_2152_elements(526)); -- 
    rr_8279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(526), ack => type_cast_3809_inst_req_0); -- 
    cr_8284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(526), ack => type_cast_3809_inst_req_1); -- 
    -- CP-element group 527:  transition  place  input  bypass 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	525 
    -- CP-element group 527: successors 
    -- CP-element group 527: 	1091 
    -- CP-element group 527:  members (5) 
      -- CP-element group 527: 	 branch_block_stmt_714/if_stmt_3799_else_link/$exit
      -- CP-element group 527: 	 branch_block_stmt_714/if_stmt_3799_else_link/else_choice_transition
      -- CP-element group 527: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1129_ifx_xthen1158
      -- CP-element group 527: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1129_ifx_xthen1158_PhiReq/$entry
      -- CP-element group 527: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1129_ifx_xthen1158_PhiReq/$exit
      -- 
    else_choice_transition_8266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 527_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3799_branch_ack_0, ack => zeropad3D_CP_2152_elements(527)); -- 
    -- CP-element group 528:  transition  input  bypass 
    -- CP-element group 528: predecessors 
    -- CP-element group 528: 	526 
    -- CP-element group 528: successors 
    -- CP-element group 528:  members (3) 
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/type_cast_3809_sample_completed_
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/type_cast_3809_Sample/$exit
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/type_cast_3809_Sample/ra
      -- 
    ra_8280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 528_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3809_inst_ack_0, ack => zeropad3D_CP_2152_elements(528)); -- 
    -- CP-element group 529:  branch  transition  place  input  output  bypass 
    -- CP-element group 529: predecessors 
    -- CP-element group 529: 	526 
    -- CP-element group 529: successors 
    -- CP-element group 529: 	530 
    -- CP-element group 529: 	531 
    -- CP-element group 529:  members (13) 
      -- CP-element group 529: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817__exit__
      -- CP-element group 529: 	 branch_block_stmt_714/if_stmt_3818__entry__
      -- CP-element group 529: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/$exit
      -- CP-element group 529: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/type_cast_3809_update_completed_
      -- CP-element group 529: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/type_cast_3809_Update/$exit
      -- CP-element group 529: 	 branch_block_stmt_714/assign_stmt_3810_to_assign_stmt_3817/type_cast_3809_Update/ca
      -- CP-element group 529: 	 branch_block_stmt_714/if_stmt_3818_dead_link/$entry
      -- CP-element group 529: 	 branch_block_stmt_714/if_stmt_3818_eval_test/$entry
      -- CP-element group 529: 	 branch_block_stmt_714/if_stmt_3818_eval_test/$exit
      -- CP-element group 529: 	 branch_block_stmt_714/if_stmt_3818_eval_test/branch_req
      -- CP-element group 529: 	 branch_block_stmt_714/R_cmp1146_3819_place
      -- CP-element group 529: 	 branch_block_stmt_714/if_stmt_3818_if_link/$entry
      -- CP-element group 529: 	 branch_block_stmt_714/if_stmt_3818_else_link/$entry
      -- 
    ca_8285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 529_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3809_inst_ack_1, ack => zeropad3D_CP_2152_elements(529)); -- 
    branch_req_8293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(529), ack => if_stmt_3818_branch_req_0); -- 
    -- CP-element group 530:  transition  place  input  bypass 
    -- CP-element group 530: predecessors 
    -- CP-element group 530: 	529 
    -- CP-element group 530: successors 
    -- CP-element group 530: 	1091 
    -- CP-element group 530:  members (5) 
      -- CP-element group 530: 	 branch_block_stmt_714/if_stmt_3818_if_link/$exit
      -- CP-element group 530: 	 branch_block_stmt_714/if_stmt_3818_if_link/if_choice_transition
      -- CP-element group 530: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1141_ifx_xthen1158
      -- CP-element group 530: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1141_ifx_xthen1158_PhiReq/$entry
      -- CP-element group 530: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1141_ifx_xthen1158_PhiReq/$exit
      -- 
    if_choice_transition_8298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 530_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3818_branch_ack_1, ack => zeropad3D_CP_2152_elements(530)); -- 
    -- CP-element group 531:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 531: predecessors 
    -- CP-element group 531: 	529 
    -- CP-element group 531: successors 
    -- CP-element group 531: 	532 
    -- CP-element group 531: 	533 
    -- CP-element group 531: 	535 
    -- CP-element group 531:  members (27) 
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843__entry__
      -- CP-element group 531: 	 branch_block_stmt_714/merge_stmt_3824__exit__
      -- CP-element group 531: 	 branch_block_stmt_714/if_stmt_3818_else_link/$exit
      -- CP-element group 531: 	 branch_block_stmt_714/if_stmt_3818_else_link/else_choice_transition
      -- CP-element group 531: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1141_lorx_xlhsx_xfalse1148
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/$entry
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_sample_start_
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_update_start_
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_word_address_calculated
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_root_address_calculated
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Sample/$entry
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Sample/word_access_start/$entry
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Sample/word_access_start/word_0/$entry
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Sample/word_access_start/word_0/rr
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Update/$entry
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Update/word_access_complete/$entry
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Update/word_access_complete/word_0/$entry
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Update/word_access_complete/word_0/cr
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/type_cast_3830_update_start_
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/type_cast_3830_Update/$entry
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/type_cast_3830_Update/cr
      -- CP-element group 531: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1141_lorx_xlhsx_xfalse1148_PhiReq/$entry
      -- CP-element group 531: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1141_lorx_xlhsx_xfalse1148_PhiReq/$exit
      -- CP-element group 531: 	 branch_block_stmt_714/merge_stmt_3824_PhiReqMerge
      -- CP-element group 531: 	 branch_block_stmt_714/merge_stmt_3824_PhiAck/$entry
      -- CP-element group 531: 	 branch_block_stmt_714/merge_stmt_3824_PhiAck/$exit
      -- CP-element group 531: 	 branch_block_stmt_714/merge_stmt_3824_PhiAck/dummy
      -- 
    else_choice_transition_8302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 531_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3818_branch_ack_0, ack => zeropad3D_CP_2152_elements(531)); -- 
    rr_8323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(531), ack => LOAD_col_high_3826_load_0_req_0); -- 
    cr_8334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(531), ack => LOAD_col_high_3826_load_0_req_1); -- 
    cr_8353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(531), ack => type_cast_3830_inst_req_1); -- 
    -- CP-element group 532:  transition  input  bypass 
    -- CP-element group 532: predecessors 
    -- CP-element group 532: 	531 
    -- CP-element group 532: successors 
    -- CP-element group 532:  members (5) 
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_sample_completed_
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Sample/$exit
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Sample/word_access_start/$exit
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Sample/word_access_start/word_0/$exit
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Sample/word_access_start/word_0/ra
      -- 
    ra_8324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 532_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3826_load_0_ack_0, ack => zeropad3D_CP_2152_elements(532)); -- 
    -- CP-element group 533:  transition  input  output  bypass 
    -- CP-element group 533: predecessors 
    -- CP-element group 533: 	531 
    -- CP-element group 533: successors 
    -- CP-element group 533: 	534 
    -- CP-element group 533:  members (12) 
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_update_completed_
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Update/$exit
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Update/word_access_complete/$exit
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Update/word_access_complete/word_0/$exit
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Update/word_access_complete/word_0/ca
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Update/LOAD_col_high_3826_Merge/$entry
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Update/LOAD_col_high_3826_Merge/$exit
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Update/LOAD_col_high_3826_Merge/merge_req
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/LOAD_col_high_3826_Update/LOAD_col_high_3826_Merge/merge_ack
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/type_cast_3830_sample_start_
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/type_cast_3830_Sample/$entry
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/type_cast_3830_Sample/rr
      -- 
    ca_8335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 533_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3826_load_0_ack_1, ack => zeropad3D_CP_2152_elements(533)); -- 
    rr_8348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(533), ack => type_cast_3830_inst_req_0); -- 
    -- CP-element group 534:  transition  input  bypass 
    -- CP-element group 534: predecessors 
    -- CP-element group 534: 	533 
    -- CP-element group 534: successors 
    -- CP-element group 534:  members (3) 
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/type_cast_3830_sample_completed_
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/type_cast_3830_Sample/$exit
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/type_cast_3830_Sample/ra
      -- 
    ra_8349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 534_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3830_inst_ack_0, ack => zeropad3D_CP_2152_elements(534)); -- 
    -- CP-element group 535:  branch  transition  place  input  output  bypass 
    -- CP-element group 535: predecessors 
    -- CP-element group 535: 	531 
    -- CP-element group 535: successors 
    -- CP-element group 535: 	536 
    -- CP-element group 535: 	537 
    -- CP-element group 535:  members (13) 
      -- CP-element group 535: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843__exit__
      -- CP-element group 535: 	 branch_block_stmt_714/if_stmt_3844__entry__
      -- CP-element group 535: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/$exit
      -- CP-element group 535: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/type_cast_3830_update_completed_
      -- CP-element group 535: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/type_cast_3830_Update/$exit
      -- CP-element group 535: 	 branch_block_stmt_714/assign_stmt_3827_to_assign_stmt_3843/type_cast_3830_Update/ca
      -- CP-element group 535: 	 branch_block_stmt_714/if_stmt_3844_dead_link/$entry
      -- CP-element group 535: 	 branch_block_stmt_714/if_stmt_3844_eval_test/$entry
      -- CP-element group 535: 	 branch_block_stmt_714/if_stmt_3844_eval_test/$exit
      -- CP-element group 535: 	 branch_block_stmt_714/if_stmt_3844_eval_test/branch_req
      -- CP-element group 535: 	 branch_block_stmt_714/R_cmp1156_3845_place
      -- CP-element group 535: 	 branch_block_stmt_714/if_stmt_3844_if_link/$entry
      -- CP-element group 535: 	 branch_block_stmt_714/if_stmt_3844_else_link/$entry
      -- 
    ca_8354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 535_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3830_inst_ack_1, ack => zeropad3D_CP_2152_elements(535)); -- 
    branch_req_8362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(535), ack => if_stmt_3844_branch_req_0); -- 
    -- CP-element group 536:  fork  transition  place  input  output  bypass 
    -- CP-element group 536: predecessors 
    -- CP-element group 536: 	535 
    -- CP-element group 536: successors 
    -- CP-element group 536: 	552 
    -- CP-element group 536: 	553 
    -- CP-element group 536: 	555 
    -- CP-element group 536: 	557 
    -- CP-element group 536: 	559 
    -- CP-element group 536: 	561 
    -- CP-element group 536: 	563 
    -- CP-element group 536: 	565 
    -- CP-element group 536: 	567 
    -- CP-element group 536: 	570 
    -- CP-element group 536:  members (46) 
      -- CP-element group 536: 	 branch_block_stmt_714/merge_stmt_3908__exit__
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013__entry__
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_update_start_
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Update/word_access_complete/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Update/word_access_complete/word_0/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/if_stmt_3844_if_link/$exit
      -- CP-element group 536: 	 branch_block_stmt_714/if_stmt_3844_if_link/if_choice_transition
      -- CP-element group 536: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1148_ifx_xelse1179
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_4008_complete/req
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_4008_complete/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3912_sample_start_
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3912_update_start_
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3912_Sample/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3912_Sample/rr
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3912_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3912_Update/cr
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3976_update_start_
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3976_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3976_Update/cr
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Update/word_access_complete/word_0/cr
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_3983_update_start_
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_final_index_sum_regn_update_start
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_final_index_sum_regn_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_final_index_sum_regn_Update/req
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_3983_complete/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_3983_complete/req
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_update_start_
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Update/word_access_complete/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Update/word_access_complete/word_0/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Update/word_access_complete/word_0/cr
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_4001_update_start_
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_4001_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_4001_Update/cr
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_4008_update_start_
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_final_index_sum_regn_update_start
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_final_index_sum_regn_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_final_index_sum_regn_Update/req
      -- CP-element group 536: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1148_ifx_xelse1179_PhiReq/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1148_ifx_xelse1179_PhiReq/$exit
      -- CP-element group 536: 	 branch_block_stmt_714/merge_stmt_3908_PhiReqMerge
      -- CP-element group 536: 	 branch_block_stmt_714/merge_stmt_3908_PhiAck/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/merge_stmt_3908_PhiAck/$exit
      -- CP-element group 536: 	 branch_block_stmt_714/merge_stmt_3908_PhiAck/dummy
      -- 
    if_choice_transition_8367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 536_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3844_branch_ack_1, ack => zeropad3D_CP_2152_elements(536)); -- 
    req_8700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(536), ack => addr_of_4008_final_reg_req_1); -- 
    rr_8525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(536), ack => type_cast_3912_inst_req_0); -- 
    cr_8530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(536), ack => type_cast_3912_inst_req_1); -- 
    cr_8544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(536), ack => type_cast_3976_inst_req_1); -- 
    cr_8750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(536), ack => ptr_deref_4011_store_0_req_1); -- 
    req_8575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(536), ack => array_obj_ref_3982_index_offset_req_1); -- 
    req_8590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(536), ack => addr_of_3983_final_reg_req_1); -- 
    cr_8635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(536), ack => ptr_deref_3987_load_0_req_1); -- 
    cr_8654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(536), ack => type_cast_4001_inst_req_1); -- 
    req_8685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(536), ack => array_obj_ref_4007_index_offset_req_1); -- 
    -- CP-element group 537:  transition  place  input  bypass 
    -- CP-element group 537: predecessors 
    -- CP-element group 537: 	535 
    -- CP-element group 537: successors 
    -- CP-element group 537: 	1091 
    -- CP-element group 537:  members (5) 
      -- CP-element group 537: 	 branch_block_stmt_714/if_stmt_3844_else_link/$exit
      -- CP-element group 537: 	 branch_block_stmt_714/if_stmt_3844_else_link/else_choice_transition
      -- CP-element group 537: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1148_ifx_xthen1158
      -- CP-element group 537: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1148_ifx_xthen1158_PhiReq/$entry
      -- CP-element group 537: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1148_ifx_xthen1158_PhiReq/$exit
      -- 
    else_choice_transition_8371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 537_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3844_branch_ack_0, ack => zeropad3D_CP_2152_elements(537)); -- 
    -- CP-element group 538:  transition  input  bypass 
    -- CP-element group 538: predecessors 
    -- CP-element group 538: 	1091 
    -- CP-element group 538: successors 
    -- CP-element group 538:  members (3) 
      -- CP-element group 538: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3854_sample_completed_
      -- CP-element group 538: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3854_Sample/$exit
      -- CP-element group 538: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3854_Sample/ra
      -- 
    ra_8385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 538_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3854_inst_ack_0, ack => zeropad3D_CP_2152_elements(538)); -- 
    -- CP-element group 539:  transition  input  bypass 
    -- CP-element group 539: predecessors 
    -- CP-element group 539: 	1091 
    -- CP-element group 539: successors 
    -- CP-element group 539: 	542 
    -- CP-element group 539:  members (3) 
      -- CP-element group 539: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3854_update_completed_
      -- CP-element group 539: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3854_Update/$exit
      -- CP-element group 539: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3854_Update/ca
      -- 
    ca_8390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 539_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3854_inst_ack_1, ack => zeropad3D_CP_2152_elements(539)); -- 
    -- CP-element group 540:  transition  input  bypass 
    -- CP-element group 540: predecessors 
    -- CP-element group 540: 	1091 
    -- CP-element group 540: successors 
    -- CP-element group 540:  members (3) 
      -- CP-element group 540: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3859_sample_completed_
      -- CP-element group 540: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3859_Sample/$exit
      -- CP-element group 540: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3859_Sample/ra
      -- 
    ra_8399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 540_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3859_inst_ack_0, ack => zeropad3D_CP_2152_elements(540)); -- 
    -- CP-element group 541:  transition  input  bypass 
    -- CP-element group 541: predecessors 
    -- CP-element group 541: 	1091 
    -- CP-element group 541: successors 
    -- CP-element group 541: 	542 
    -- CP-element group 541:  members (3) 
      -- CP-element group 541: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3859_update_completed_
      -- CP-element group 541: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3859_Update/$exit
      -- CP-element group 541: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3859_Update/ca
      -- 
    ca_8404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 541_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3859_inst_ack_1, ack => zeropad3D_CP_2152_elements(541)); -- 
    -- CP-element group 542:  join  transition  output  bypass 
    -- CP-element group 542: predecessors 
    -- CP-element group 542: 	539 
    -- CP-element group 542: 	541 
    -- CP-element group 542: successors 
    -- CP-element group 542: 	543 
    -- CP-element group 542:  members (3) 
      -- CP-element group 542: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3893_sample_start_
      -- CP-element group 542: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3893_Sample/$entry
      -- CP-element group 542: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3893_Sample/rr
      -- 
    rr_8412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(542), ack => type_cast_3893_inst_req_0); -- 
    zeropad3D_cp_element_group_542: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_542"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(539) & zeropad3D_CP_2152_elements(541);
      gj_zeropad3D_cp_element_group_542 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(542), clk => clk, reset => reset); --
    end block;
    -- CP-element group 543:  transition  input  bypass 
    -- CP-element group 543: predecessors 
    -- CP-element group 543: 	542 
    -- CP-element group 543: successors 
    -- CP-element group 543:  members (3) 
      -- CP-element group 543: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3893_sample_completed_
      -- CP-element group 543: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3893_Sample/$exit
      -- CP-element group 543: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3893_Sample/ra
      -- 
    ra_8413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 543_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3893_inst_ack_0, ack => zeropad3D_CP_2152_elements(543)); -- 
    -- CP-element group 544:  transition  input  output  bypass 
    -- CP-element group 544: predecessors 
    -- CP-element group 544: 	1091 
    -- CP-element group 544: successors 
    -- CP-element group 544: 	545 
    -- CP-element group 544:  members (16) 
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3893_update_completed_
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3893_Update/$exit
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3893_Update/ca
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_index_resized_1
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_index_scaled_1
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_index_computed_1
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_index_resize_1/$entry
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_index_resize_1/$exit
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_index_resize_1/index_resize_req
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_index_resize_1/index_resize_ack
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_index_scale_1/$entry
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_index_scale_1/$exit
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_index_scale_1/scale_rename_req
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_index_scale_1/scale_rename_ack
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_final_index_sum_regn_Sample/$entry
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_final_index_sum_regn_Sample/req
      -- 
    ca_8418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 544_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3893_inst_ack_1, ack => zeropad3D_CP_2152_elements(544)); -- 
    req_8443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(544), ack => array_obj_ref_3899_index_offset_req_0); -- 
    -- CP-element group 545:  transition  input  bypass 
    -- CP-element group 545: predecessors 
    -- CP-element group 545: 	544 
    -- CP-element group 545: successors 
    -- CP-element group 545: 	551 
    -- CP-element group 545:  members (3) 
      -- CP-element group 545: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_final_index_sum_regn_sample_complete
      -- CP-element group 545: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_final_index_sum_regn_Sample/$exit
      -- CP-element group 545: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_final_index_sum_regn_Sample/ack
      -- 
    ack_8444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 545_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3899_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(545)); -- 
    -- CP-element group 546:  transition  input  output  bypass 
    -- CP-element group 546: predecessors 
    -- CP-element group 546: 	1091 
    -- CP-element group 546: successors 
    -- CP-element group 546: 	547 
    -- CP-element group 546:  members (11) 
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/addr_of_3900_sample_start_
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_root_address_calculated
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_offset_calculated
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_final_index_sum_regn_Update/$exit
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_final_index_sum_regn_Update/ack
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_base_plus_offset/$entry
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_base_plus_offset/$exit
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_base_plus_offset/sum_rename_req
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_base_plus_offset/sum_rename_ack
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/addr_of_3900_request/$entry
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/addr_of_3900_request/req
      -- 
    ack_8449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 546_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3899_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(546)); -- 
    req_8458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(546), ack => addr_of_3900_final_reg_req_0); -- 
    -- CP-element group 547:  transition  input  bypass 
    -- CP-element group 547: predecessors 
    -- CP-element group 547: 	546 
    -- CP-element group 547: successors 
    -- CP-element group 547:  members (3) 
      -- CP-element group 547: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/addr_of_3900_sample_completed_
      -- CP-element group 547: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/addr_of_3900_request/$exit
      -- CP-element group 547: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/addr_of_3900_request/ack
      -- 
    ack_8459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 547_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3900_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(547)); -- 
    -- CP-element group 548:  join  fork  transition  input  output  bypass 
    -- CP-element group 548: predecessors 
    -- CP-element group 548: 	1091 
    -- CP-element group 548: successors 
    -- CP-element group 548: 	549 
    -- CP-element group 548:  members (28) 
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/addr_of_3900_update_completed_
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/addr_of_3900_complete/$exit
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/addr_of_3900_complete/ack
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_sample_start_
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_base_address_calculated
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_word_address_calculated
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_root_address_calculated
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_base_address_resized
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_base_addr_resize/$entry
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_base_addr_resize/$exit
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_base_addr_resize/base_resize_req
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_base_addr_resize/base_resize_ack
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_base_plus_offset/$entry
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_base_plus_offset/$exit
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_base_plus_offset/sum_rename_req
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_base_plus_offset/sum_rename_ack
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_word_addrgen/$entry
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_word_addrgen/$exit
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_word_addrgen/root_register_req
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_word_addrgen/root_register_ack
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Sample/$entry
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Sample/ptr_deref_3903_Split/$entry
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Sample/ptr_deref_3903_Split/$exit
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Sample/ptr_deref_3903_Split/split_req
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Sample/ptr_deref_3903_Split/split_ack
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Sample/word_access_start/$entry
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Sample/word_access_start/word_0/$entry
      -- CP-element group 548: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Sample/word_access_start/word_0/rr
      -- 
    ack_8464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 548_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3900_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(548)); -- 
    rr_8502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(548), ack => ptr_deref_3903_store_0_req_0); -- 
    -- CP-element group 549:  transition  input  bypass 
    -- CP-element group 549: predecessors 
    -- CP-element group 549: 	548 
    -- CP-element group 549: successors 
    -- CP-element group 549:  members (5) 
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_sample_completed_
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Sample/$exit
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Sample/word_access_start/$exit
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Sample/word_access_start/word_0/$exit
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Sample/word_access_start/word_0/ra
      -- 
    ra_8503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 549_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3903_store_0_ack_0, ack => zeropad3D_CP_2152_elements(549)); -- 
    -- CP-element group 550:  transition  input  bypass 
    -- CP-element group 550: predecessors 
    -- CP-element group 550: 	1091 
    -- CP-element group 550: successors 
    -- CP-element group 550: 	551 
    -- CP-element group 550:  members (5) 
      -- CP-element group 550: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_update_completed_
      -- CP-element group 550: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Update/$exit
      -- CP-element group 550: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Update/word_access_complete/$exit
      -- CP-element group 550: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Update/word_access_complete/word_0/$exit
      -- CP-element group 550: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Update/word_access_complete/word_0/ca
      -- 
    ca_8514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 550_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3903_store_0_ack_1, ack => zeropad3D_CP_2152_elements(550)); -- 
    -- CP-element group 551:  join  transition  place  bypass 
    -- CP-element group 551: predecessors 
    -- CP-element group 551: 	545 
    -- CP-element group 551: 	550 
    -- CP-element group 551: successors 
    -- CP-element group 551: 	1092 
    -- CP-element group 551:  members (5) 
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906__exit__
      -- CP-element group 551: 	 branch_block_stmt_714/ifx_xthen1158_ifx_xend1227
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/$exit
      -- CP-element group 551: 	 branch_block_stmt_714/ifx_xthen1158_ifx_xend1227_PhiReq/$entry
      -- CP-element group 551: 	 branch_block_stmt_714/ifx_xthen1158_ifx_xend1227_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_551: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_551"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(545) & zeropad3D_CP_2152_elements(550);
      gj_zeropad3D_cp_element_group_551 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(551), clk => clk, reset => reset); --
    end block;
    -- CP-element group 552:  transition  input  bypass 
    -- CP-element group 552: predecessors 
    -- CP-element group 552: 	536 
    -- CP-element group 552: successors 
    -- CP-element group 552:  members (3) 
      -- CP-element group 552: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3912_sample_completed_
      -- CP-element group 552: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3912_Sample/$exit
      -- CP-element group 552: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3912_Sample/ra
      -- 
    ra_8526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 552_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3912_inst_ack_0, ack => zeropad3D_CP_2152_elements(552)); -- 
    -- CP-element group 553:  fork  transition  input  output  bypass 
    -- CP-element group 553: predecessors 
    -- CP-element group 553: 	536 
    -- CP-element group 553: successors 
    -- CP-element group 553: 	554 
    -- CP-element group 553: 	562 
    -- CP-element group 553:  members (9) 
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3912_update_completed_
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3912_Update/$exit
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3912_Update/ca
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3976_sample_start_
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3976_Sample/$entry
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3976_Sample/rr
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_4001_sample_start_
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_4001_Sample/$entry
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_4001_Sample/rr
      -- 
    ca_8531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 553_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3912_inst_ack_1, ack => zeropad3D_CP_2152_elements(553)); -- 
    rr_8539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(553), ack => type_cast_3976_inst_req_0); -- 
    rr_8649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(553), ack => type_cast_4001_inst_req_0); -- 
    -- CP-element group 554:  transition  input  bypass 
    -- CP-element group 554: predecessors 
    -- CP-element group 554: 	553 
    -- CP-element group 554: successors 
    -- CP-element group 554:  members (3) 
      -- CP-element group 554: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3976_sample_completed_
      -- CP-element group 554: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3976_Sample/$exit
      -- CP-element group 554: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3976_Sample/ra
      -- 
    ra_8540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 554_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3976_inst_ack_0, ack => zeropad3D_CP_2152_elements(554)); -- 
    -- CP-element group 555:  transition  input  output  bypass 
    -- CP-element group 555: predecessors 
    -- CP-element group 555: 	536 
    -- CP-element group 555: successors 
    -- CP-element group 555: 	556 
    -- CP-element group 555:  members (16) 
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3976_update_completed_
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3976_Update/$exit
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_3976_Update/ca
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_index_resized_1
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_index_scaled_1
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_index_computed_1
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_index_resize_1/$entry
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_index_resize_1/$exit
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_index_resize_1/index_resize_req
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_index_resize_1/index_resize_ack
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_index_scale_1/$entry
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_index_scale_1/$exit
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_index_scale_1/scale_rename_req
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_index_scale_1/scale_rename_ack
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_final_index_sum_regn_Sample/$entry
      -- CP-element group 555: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_final_index_sum_regn_Sample/req
      -- 
    ca_8545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 555_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3976_inst_ack_1, ack => zeropad3D_CP_2152_elements(555)); -- 
    req_8570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(555), ack => array_obj_ref_3982_index_offset_req_0); -- 
    -- CP-element group 556:  transition  input  bypass 
    -- CP-element group 556: predecessors 
    -- CP-element group 556: 	555 
    -- CP-element group 556: successors 
    -- CP-element group 556: 	571 
    -- CP-element group 556:  members (3) 
      -- CP-element group 556: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_final_index_sum_regn_sample_complete
      -- CP-element group 556: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_final_index_sum_regn_Sample/$exit
      -- CP-element group 556: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_final_index_sum_regn_Sample/ack
      -- 
    ack_8571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 556_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3982_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(556)); -- 
    -- CP-element group 557:  transition  input  output  bypass 
    -- CP-element group 557: predecessors 
    -- CP-element group 557: 	536 
    -- CP-element group 557: successors 
    -- CP-element group 557: 	558 
    -- CP-element group 557:  members (11) 
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_3983_sample_start_
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_root_address_calculated
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_offset_calculated
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_final_index_sum_regn_Update/$exit
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_final_index_sum_regn_Update/ack
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_base_plus_offset/$entry
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_base_plus_offset/$exit
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_base_plus_offset/sum_rename_req
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_3982_base_plus_offset/sum_rename_ack
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_3983_request/$entry
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_3983_request/req
      -- 
    ack_8576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 557_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3982_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(557)); -- 
    req_8585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(557), ack => addr_of_3983_final_reg_req_0); -- 
    -- CP-element group 558:  transition  input  bypass 
    -- CP-element group 558: predecessors 
    -- CP-element group 558: 	557 
    -- CP-element group 558: successors 
    -- CP-element group 558:  members (3) 
      -- CP-element group 558: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_3983_sample_completed_
      -- CP-element group 558: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_3983_request/$exit
      -- CP-element group 558: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_3983_request/ack
      -- 
    ack_8586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 558_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3983_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(558)); -- 
    -- CP-element group 559:  join  fork  transition  input  output  bypass 
    -- CP-element group 559: predecessors 
    -- CP-element group 559: 	536 
    -- CP-element group 559: successors 
    -- CP-element group 559: 	560 
    -- CP-element group 559:  members (24) 
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_3983_update_completed_
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_3983_complete/$exit
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_3983_complete/ack
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_sample_start_
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_base_address_calculated
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_word_address_calculated
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_root_address_calculated
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_base_address_resized
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_base_addr_resize/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_base_addr_resize/$exit
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_base_addr_resize/base_resize_req
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_base_addr_resize/base_resize_ack
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_base_plus_offset/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_base_plus_offset/$exit
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_base_plus_offset/sum_rename_req
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_base_plus_offset/sum_rename_ack
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_word_addrgen/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_word_addrgen/$exit
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_word_addrgen/root_register_req
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_word_addrgen/root_register_ack
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Sample/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Sample/word_access_start/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Sample/word_access_start/word_0/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Sample/word_access_start/word_0/rr
      -- 
    ack_8591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 559_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3983_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(559)); -- 
    rr_8624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(559), ack => ptr_deref_3987_load_0_req_0); -- 
    -- CP-element group 560:  transition  input  bypass 
    -- CP-element group 560: predecessors 
    -- CP-element group 560: 	559 
    -- CP-element group 560: successors 
    -- CP-element group 560:  members (5) 
      -- CP-element group 560: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_sample_completed_
      -- CP-element group 560: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Sample/$exit
      -- CP-element group 560: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Sample/word_access_start/$exit
      -- CP-element group 560: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Sample/word_access_start/word_0/$exit
      -- CP-element group 560: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Sample/word_access_start/word_0/ra
      -- 
    ra_8625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 560_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3987_load_0_ack_0, ack => zeropad3D_CP_2152_elements(560)); -- 
    -- CP-element group 561:  transition  input  bypass 
    -- CP-element group 561: predecessors 
    -- CP-element group 561: 	536 
    -- CP-element group 561: successors 
    -- CP-element group 561: 	568 
    -- CP-element group 561:  members (9) 
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_update_completed_
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Update/$exit
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Update/word_access_complete/$exit
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Update/word_access_complete/word_0/$exit
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Update/word_access_complete/word_0/ca
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Update/ptr_deref_3987_Merge/$entry
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Update/ptr_deref_3987_Merge/$exit
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Update/ptr_deref_3987_Merge/merge_req
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_3987_Update/ptr_deref_3987_Merge/merge_ack
      -- 
    ca_8636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 561_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3987_load_0_ack_1, ack => zeropad3D_CP_2152_elements(561)); -- 
    -- CP-element group 562:  transition  input  bypass 
    -- CP-element group 562: predecessors 
    -- CP-element group 562: 	553 
    -- CP-element group 562: successors 
    -- CP-element group 562:  members (3) 
      -- CP-element group 562: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_4001_sample_completed_
      -- CP-element group 562: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_4001_Sample/$exit
      -- CP-element group 562: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_4001_Sample/ra
      -- 
    ra_8650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 562_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4001_inst_ack_0, ack => zeropad3D_CP_2152_elements(562)); -- 
    -- CP-element group 563:  transition  input  output  bypass 
    -- CP-element group 563: predecessors 
    -- CP-element group 563: 	536 
    -- CP-element group 563: successors 
    -- CP-element group 563: 	564 
    -- CP-element group 563:  members (16) 
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_4001_update_completed_
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_4001_Update/$exit
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/type_cast_4001_Update/ca
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_index_resized_1
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_index_scaled_1
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_index_computed_1
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_index_resize_1/$entry
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_index_resize_1/$exit
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_index_resize_1/index_resize_req
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_index_resize_1/index_resize_ack
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_index_scale_1/$entry
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_index_scale_1/$exit
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_index_scale_1/scale_rename_req
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_index_scale_1/scale_rename_ack
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_final_index_sum_regn_Sample/$entry
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_final_index_sum_regn_Sample/req
      -- 
    ca_8655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 563_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4001_inst_ack_1, ack => zeropad3D_CP_2152_elements(563)); -- 
    req_8680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(563), ack => array_obj_ref_4007_index_offset_req_0); -- 
    -- CP-element group 564:  transition  input  bypass 
    -- CP-element group 564: predecessors 
    -- CP-element group 564: 	563 
    -- CP-element group 564: successors 
    -- CP-element group 564: 	571 
    -- CP-element group 564:  members (3) 
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_final_index_sum_regn_sample_complete
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_final_index_sum_regn_Sample/$exit
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_final_index_sum_regn_Sample/ack
      -- 
    ack_8681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 564_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4007_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(564)); -- 
    -- CP-element group 565:  transition  input  output  bypass 
    -- CP-element group 565: predecessors 
    -- CP-element group 565: 	536 
    -- CP-element group 565: successors 
    -- CP-element group 565: 	566 
    -- CP-element group 565:  members (11) 
      -- CP-element group 565: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_4008_request/req
      -- CP-element group 565: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_4008_request/$entry
      -- CP-element group 565: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_4008_sample_start_
      -- CP-element group 565: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_root_address_calculated
      -- CP-element group 565: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_offset_calculated
      -- CP-element group 565: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_final_index_sum_regn_Update/$exit
      -- CP-element group 565: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_final_index_sum_regn_Update/ack
      -- CP-element group 565: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_base_plus_offset/$entry
      -- CP-element group 565: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_base_plus_offset/$exit
      -- CP-element group 565: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_base_plus_offset/sum_rename_req
      -- CP-element group 565: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/array_obj_ref_4007_base_plus_offset/sum_rename_ack
      -- 
    ack_8686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 565_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4007_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(565)); -- 
    req_8695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(565), ack => addr_of_4008_final_reg_req_0); -- 
    -- CP-element group 566:  transition  input  bypass 
    -- CP-element group 566: predecessors 
    -- CP-element group 566: 	565 
    -- CP-element group 566: successors 
    -- CP-element group 566:  members (3) 
      -- CP-element group 566: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_4008_request/ack
      -- CP-element group 566: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_4008_request/$exit
      -- CP-element group 566: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_4008_sample_completed_
      -- 
    ack_8696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 566_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4008_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(566)); -- 
    -- CP-element group 567:  fork  transition  input  bypass 
    -- CP-element group 567: predecessors 
    -- CP-element group 567: 	536 
    -- CP-element group 567: successors 
    -- CP-element group 567: 	568 
    -- CP-element group 567:  members (19) 
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_base_address_calculated
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_word_address_calculated
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_root_address_calculated
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_base_address_resized
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_base_addr_resize/$entry
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_base_addr_resize/$exit
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_base_addr_resize/base_resize_req
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_base_addr_resize/base_resize_ack
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_word_addrgen/root_register_ack
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_word_addrgen/root_register_req
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_word_addrgen/$exit
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_word_addrgen/$entry
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_base_plus_offset/sum_rename_ack
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_base_plus_offset/sum_rename_req
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_base_plus_offset/$exit
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_base_plus_offset/$entry
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_4008_complete/ack
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_4008_complete/$exit
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/addr_of_4008_update_completed_
      -- 
    ack_8701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 567_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4008_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(567)); -- 
    -- CP-element group 568:  join  transition  output  bypass 
    -- CP-element group 568: predecessors 
    -- CP-element group 568: 	561 
    -- CP-element group 568: 	567 
    -- CP-element group 568: successors 
    -- CP-element group 568: 	569 
    -- CP-element group 568:  members (9) 
      -- CP-element group 568: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Sample/word_access_start/word_0/rr
      -- CP-element group 568: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Sample/word_access_start/word_0/$entry
      -- CP-element group 568: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Sample/word_access_start/$entry
      -- CP-element group 568: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Sample/ptr_deref_4011_Split/split_ack
      -- CP-element group 568: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Sample/ptr_deref_4011_Split/split_req
      -- CP-element group 568: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Sample/ptr_deref_4011_Split/$exit
      -- CP-element group 568: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Sample/ptr_deref_4011_Split/$entry
      -- CP-element group 568: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Sample/$entry
      -- CP-element group 568: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_sample_start_
      -- 
    rr_8739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(568), ack => ptr_deref_4011_store_0_req_0); -- 
    zeropad3D_cp_element_group_568: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_568"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(561) & zeropad3D_CP_2152_elements(567);
      gj_zeropad3D_cp_element_group_568 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(568), clk => clk, reset => reset); --
    end block;
    -- CP-element group 569:  transition  input  bypass 
    -- CP-element group 569: predecessors 
    -- CP-element group 569: 	568 
    -- CP-element group 569: successors 
    -- CP-element group 569:  members (5) 
      -- CP-element group 569: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Sample/word_access_start/word_0/ra
      -- CP-element group 569: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Sample/word_access_start/word_0/$exit
      -- CP-element group 569: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Sample/word_access_start/$exit
      -- CP-element group 569: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_sample_completed_
      -- CP-element group 569: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Sample/$exit
      -- 
    ra_8740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 569_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4011_store_0_ack_0, ack => zeropad3D_CP_2152_elements(569)); -- 
    -- CP-element group 570:  transition  input  bypass 
    -- CP-element group 570: predecessors 
    -- CP-element group 570: 	536 
    -- CP-element group 570: successors 
    -- CP-element group 570: 	571 
    -- CP-element group 570:  members (5) 
      -- CP-element group 570: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Update/$exit
      -- CP-element group 570: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_update_completed_
      -- CP-element group 570: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Update/word_access_complete/$exit
      -- CP-element group 570: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Update/word_access_complete/word_0/ca
      -- CP-element group 570: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/ptr_deref_4011_Update/word_access_complete/word_0/$exit
      -- 
    ca_8751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 570_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4011_store_0_ack_1, ack => zeropad3D_CP_2152_elements(570)); -- 
    -- CP-element group 571:  join  transition  place  bypass 
    -- CP-element group 571: predecessors 
    -- CP-element group 571: 	556 
    -- CP-element group 571: 	564 
    -- CP-element group 571: 	570 
    -- CP-element group 571: successors 
    -- CP-element group 571: 	1092 
    -- CP-element group 571:  members (5) 
      -- CP-element group 571: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013__exit__
      -- CP-element group 571: 	 branch_block_stmt_714/ifx_xelse1179_ifx_xend1227
      -- CP-element group 571: 	 branch_block_stmt_714/assign_stmt_3913_to_assign_stmt_4013/$exit
      -- CP-element group 571: 	 branch_block_stmt_714/ifx_xelse1179_ifx_xend1227_PhiReq/$entry
      -- CP-element group 571: 	 branch_block_stmt_714/ifx_xelse1179_ifx_xend1227_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_571: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_571"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(556) & zeropad3D_CP_2152_elements(564) & zeropad3D_CP_2152_elements(570);
      gj_zeropad3D_cp_element_group_571 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(571), clk => clk, reset => reset); --
    end block;
    -- CP-element group 572:  transition  input  bypass 
    -- CP-element group 572: predecessors 
    -- CP-element group 572: 	1092 
    -- CP-element group 572: successors 
    -- CP-element group 572:  members (3) 
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/type_cast_4019_Sample/ra
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/type_cast_4019_Sample/$exit
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/type_cast_4019_sample_completed_
      -- 
    ra_8763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 572_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4019_inst_ack_0, ack => zeropad3D_CP_2152_elements(572)); -- 
    -- CP-element group 573:  branch  transition  place  input  output  bypass 
    -- CP-element group 573: predecessors 
    -- CP-element group 573: 	1092 
    -- CP-element group 573: successors 
    -- CP-element group 573: 	574 
    -- CP-element group 573: 	575 
    -- CP-element group 573:  members (13) 
      -- CP-element group 573: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033__exit__
      -- CP-element group 573: 	 branch_block_stmt_714/if_stmt_4034__entry__
      -- CP-element group 573: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/type_cast_4019_Update/$exit
      -- CP-element group 573: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/type_cast_4019_Update/ca
      -- CP-element group 573: 	 branch_block_stmt_714/if_stmt_4034_dead_link/$entry
      -- CP-element group 573: 	 branch_block_stmt_714/if_stmt_4034_eval_test/$entry
      -- CP-element group 573: 	 branch_block_stmt_714/if_stmt_4034_eval_test/$exit
      -- CP-element group 573: 	 branch_block_stmt_714/if_stmt_4034_eval_test/branch_req
      -- CP-element group 573: 	 branch_block_stmt_714/if_stmt_4034_if_link/$entry
      -- CP-element group 573: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/type_cast_4019_update_completed_
      -- CP-element group 573: 	 branch_block_stmt_714/if_stmt_4034_else_link/$entry
      -- CP-element group 573: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/$exit
      -- CP-element group 573: 	 branch_block_stmt_714/R_cmp1235_4035_place
      -- 
    ca_8768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 573_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4019_inst_ack_1, ack => zeropad3D_CP_2152_elements(573)); -- 
    branch_req_8776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(573), ack => if_stmt_4034_branch_req_0); -- 
    -- CP-element group 574:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 574: predecessors 
    -- CP-element group 574: 	573 
    -- CP-element group 574: successors 
    -- CP-element group 574: 	1101 
    -- CP-element group 574: 	1102 
    -- CP-element group 574: 	1104 
    -- CP-element group 574: 	1105 
    -- CP-element group 574: 	1107 
    -- CP-element group 574: 	1108 
    -- CP-element group 574:  members (40) 
      -- CP-element group 574: 	 branch_block_stmt_714/merge_stmt_4040__exit__
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_4046__entry__
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_4046__exit__
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_4046/$exit
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_4046/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xend1227_ifx_xthen1237
      -- CP-element group 574: 	 branch_block_stmt_714/if_stmt_4034_if_link/if_choice_transition
      -- CP-element group 574: 	 branch_block_stmt_714/if_stmt_4034_if_link/$exit
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xend1227_ifx_xthen1237_PhiReq/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xend1227_ifx_xthen1237_PhiReq/$exit
      -- CP-element group 574: 	 branch_block_stmt_714/merge_stmt_4040_PhiReqMerge
      -- CP-element group 574: 	 branch_block_stmt_714/merge_stmt_4040_PhiAck/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/merge_stmt_4040_PhiAck/$exit
      -- CP-element group 574: 	 branch_block_stmt_714/merge_stmt_4040_PhiAck/dummy
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/type_cast_4136/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/type_cast_4136/SplitProtocol/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/type_cast_4136/SplitProtocol/Sample/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/type_cast_4136/SplitProtocol/Sample/rr
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/type_cast_4136/SplitProtocol/Update/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/type_cast_4136/SplitProtocol/Update/cr
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4143/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4143/SplitProtocol/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4143/SplitProtocol/Sample/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4143/SplitProtocol/Sample/rr
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4143/SplitProtocol/Update/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4143/SplitProtocol/Update/cr
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4149/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4149/SplitProtocol/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4149/SplitProtocol/Sample/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4149/SplitProtocol/Sample/rr
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4149/SplitProtocol/Update/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4149/SplitProtocol/Update/cr
      -- 
    if_choice_transition_8781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 574_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4034_branch_ack_1, ack => zeropad3D_CP_2152_elements(574)); -- 
    rr_13391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(574), ack => type_cast_4136_inst_req_0); -- 
    cr_13396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(574), ack => type_cast_4136_inst_req_1); -- 
    rr_13414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(574), ack => type_cast_4143_inst_req_0); -- 
    cr_13419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(574), ack => type_cast_4143_inst_req_1); -- 
    rr_13437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(574), ack => type_cast_4149_inst_req_0); -- 
    cr_13442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(574), ack => type_cast_4149_inst_req_1); -- 
    -- CP-element group 575:  fork  transition  place  input  output  bypass 
    -- CP-element group 575: predecessors 
    -- CP-element group 575: 	573 
    -- CP-element group 575: successors 
    -- CP-element group 575: 	576 
    -- CP-element group 575: 	577 
    -- CP-element group 575: 	578 
    -- CP-element group 575: 	579 
    -- CP-element group 575: 	581 
    -- CP-element group 575: 	584 
    -- CP-element group 575: 	586 
    -- CP-element group 575: 	587 
    -- CP-element group 575: 	588 
    -- CP-element group 575: 	590 
    -- CP-element group 575:  members (54) 
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125__entry__
      -- CP-element group 575: 	 branch_block_stmt_714/merge_stmt_4048__exit__
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4095_Update/cr
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_sample_start_
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4065_Update/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4065_Update/cr
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_update_start_
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4058_sample_start_
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_word_address_calculated
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4102_Update/cr
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4095_Update/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4102_Update/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4065_update_start_
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4095_update_start_
      -- CP-element group 575: 	 branch_block_stmt_714/if_stmt_4034_else_link/else_choice_transition
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4079_Update/cr
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Update/word_access_complete/word_0/cr
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4079_Update/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/if_stmt_4034_else_link/$exit
      -- CP-element group 575: 	 branch_block_stmt_714/ifx_xend1227_ifx_xelse1242
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4102_update_start_
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Update/word_access_complete/word_0/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Update/word_access_complete/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Update/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Update/word_access_complete/word_0/cr
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Sample/word_access_start/word_0/rr
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Update/word_access_complete/word_0/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Update/word_access_complete/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Sample/word_access_start/word_0/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Update/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Sample/word_access_start/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Sample/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Sample/word_access_start/word_0/rr
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_root_address_calculated
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_word_address_calculated
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Sample/word_access_start/word_0/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_update_start_
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4079_update_start_
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Sample/word_access_start/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_sample_start_
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Sample/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_root_address_calculated
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4058_Update/cr
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4058_Update/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4058_Sample/rr
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4058_Sample/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4058_update_start_
      -- CP-element group 575: 	 branch_block_stmt_714/ifx_xend1227_ifx_xelse1242_PhiReq/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/ifx_xend1227_ifx_xelse1242_PhiReq/$exit
      -- CP-element group 575: 	 branch_block_stmt_714/merge_stmt_4048_PhiReqMerge
      -- CP-element group 575: 	 branch_block_stmt_714/merge_stmt_4048_PhiAck/$entry
      -- CP-element group 575: 	 branch_block_stmt_714/merge_stmt_4048_PhiAck/$exit
      -- CP-element group 575: 	 branch_block_stmt_714/merge_stmt_4048_PhiAck/dummy
      -- 
    else_choice_transition_8785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 575_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4034_branch_ack_0, ack => zeropad3D_CP_2152_elements(575)); -- 
    cr_8881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(575), ack => type_cast_4095_inst_req_1); -- 
    cr_8853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(575), ack => type_cast_4065_inst_req_1); -- 
    cr_8928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(575), ack => type_cast_4102_inst_req_1); -- 
    cr_8867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(575), ack => type_cast_4079_inst_req_1); -- 
    cr_8834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(575), ack => LOAD_col_high_4061_load_0_req_1); -- 
    cr_8909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(575), ack => LOAD_row_high_4098_load_0_req_1); -- 
    rr_8823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(575), ack => LOAD_col_high_4061_load_0_req_0); -- 
    rr_8898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(575), ack => LOAD_row_high_4098_load_0_req_0); -- 
    cr_8806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(575), ack => type_cast_4058_inst_req_1); -- 
    rr_8801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(575), ack => type_cast_4058_inst_req_0); -- 
    -- CP-element group 576:  transition  input  bypass 
    -- CP-element group 576: predecessors 
    -- CP-element group 576: 	575 
    -- CP-element group 576: successors 
    -- CP-element group 576:  members (3) 
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4058_sample_completed_
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4058_Sample/ra
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4058_Sample/$exit
      -- 
    ra_8802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 576_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4058_inst_ack_0, ack => zeropad3D_CP_2152_elements(576)); -- 
    -- CP-element group 577:  transition  input  bypass 
    -- CP-element group 577: predecessors 
    -- CP-element group 577: 	575 
    -- CP-element group 577: successors 
    -- CP-element group 577: 	582 
    -- CP-element group 577:  members (3) 
      -- CP-element group 577: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4058_Update/ca
      -- CP-element group 577: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4058_Update/$exit
      -- CP-element group 577: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4058_update_completed_
      -- 
    ca_8807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 577_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4058_inst_ack_1, ack => zeropad3D_CP_2152_elements(577)); -- 
    -- CP-element group 578:  transition  input  bypass 
    -- CP-element group 578: predecessors 
    -- CP-element group 578: 	575 
    -- CP-element group 578: successors 
    -- CP-element group 578:  members (5) 
      -- CP-element group 578: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Sample/word_access_start/word_0/ra
      -- CP-element group 578: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Sample/word_access_start/word_0/$exit
      -- CP-element group 578: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Sample/word_access_start/$exit
      -- CP-element group 578: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Sample/$exit
      -- CP-element group 578: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_sample_completed_
      -- 
    ra_8824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 578_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4061_load_0_ack_0, ack => zeropad3D_CP_2152_elements(578)); -- 
    -- CP-element group 579:  transition  input  output  bypass 
    -- CP-element group 579: predecessors 
    -- CP-element group 579: 	575 
    -- CP-element group 579: successors 
    -- CP-element group 579: 	580 
    -- CP-element group 579:  members (12) 
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4065_Sample/rr
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4065_Sample/$entry
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4065_sample_start_
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Update/LOAD_col_high_4061_Merge/merge_ack
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Update/LOAD_col_high_4061_Merge/merge_req
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Update/LOAD_col_high_4061_Merge/$exit
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Update/LOAD_col_high_4061_Merge/$entry
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Update/word_access_complete/word_0/ca
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Update/word_access_complete/word_0/$exit
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Update/word_access_complete/$exit
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_Update/$exit
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_col_high_4061_update_completed_
      -- 
    ca_8835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 579_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4061_load_0_ack_1, ack => zeropad3D_CP_2152_elements(579)); -- 
    rr_8848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(579), ack => type_cast_4065_inst_req_0); -- 
    -- CP-element group 580:  transition  input  bypass 
    -- CP-element group 580: predecessors 
    -- CP-element group 580: 	579 
    -- CP-element group 580: successors 
    -- CP-element group 580:  members (3) 
      -- CP-element group 580: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4065_Sample/ra
      -- CP-element group 580: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4065_Sample/$exit
      -- CP-element group 580: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4065_sample_completed_
      -- 
    ra_8849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 580_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4065_inst_ack_0, ack => zeropad3D_CP_2152_elements(580)); -- 
    -- CP-element group 581:  transition  input  bypass 
    -- CP-element group 581: predecessors 
    -- CP-element group 581: 	575 
    -- CP-element group 581: successors 
    -- CP-element group 581: 	582 
    -- CP-element group 581:  members (3) 
      -- CP-element group 581: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4065_Update/$exit
      -- CP-element group 581: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4065_Update/ca
      -- CP-element group 581: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4065_update_completed_
      -- 
    ca_8854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 581_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4065_inst_ack_1, ack => zeropad3D_CP_2152_elements(581)); -- 
    -- CP-element group 582:  join  transition  output  bypass 
    -- CP-element group 582: predecessors 
    -- CP-element group 582: 	577 
    -- CP-element group 582: 	581 
    -- CP-element group 582: successors 
    -- CP-element group 582: 	583 
    -- CP-element group 582:  members (3) 
      -- CP-element group 582: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4079_sample_start_
      -- CP-element group 582: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4079_Sample/rr
      -- CP-element group 582: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4079_Sample/$entry
      -- 
    rr_8862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(582), ack => type_cast_4079_inst_req_0); -- 
    zeropad3D_cp_element_group_582: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_582"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(577) & zeropad3D_CP_2152_elements(581);
      gj_zeropad3D_cp_element_group_582 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(582), clk => clk, reset => reset); --
    end block;
    -- CP-element group 583:  transition  input  bypass 
    -- CP-element group 583: predecessors 
    -- CP-element group 583: 	582 
    -- CP-element group 583: successors 
    -- CP-element group 583:  members (3) 
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4079_sample_completed_
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4079_Sample/ra
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4079_Sample/$exit
      -- 
    ra_8863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 583_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4079_inst_ack_0, ack => zeropad3D_CP_2152_elements(583)); -- 
    -- CP-element group 584:  transition  input  output  bypass 
    -- CP-element group 584: predecessors 
    -- CP-element group 584: 	575 
    -- CP-element group 584: successors 
    -- CP-element group 584: 	585 
    -- CP-element group 584:  members (6) 
      -- CP-element group 584: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4095_Sample/rr
      -- CP-element group 584: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4095_Sample/$entry
      -- CP-element group 584: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4095_sample_start_
      -- CP-element group 584: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4079_Update/ca
      -- CP-element group 584: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4079_Update/$exit
      -- CP-element group 584: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4079_update_completed_
      -- 
    ca_8868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 584_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4079_inst_ack_1, ack => zeropad3D_CP_2152_elements(584)); -- 
    rr_8876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(584), ack => type_cast_4095_inst_req_0); -- 
    -- CP-element group 585:  transition  input  bypass 
    -- CP-element group 585: predecessors 
    -- CP-element group 585: 	584 
    -- CP-element group 585: successors 
    -- CP-element group 585:  members (3) 
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4095_Sample/ra
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4095_Sample/$exit
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4095_sample_completed_
      -- 
    ra_8877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 585_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4095_inst_ack_0, ack => zeropad3D_CP_2152_elements(585)); -- 
    -- CP-element group 586:  transition  input  bypass 
    -- CP-element group 586: predecessors 
    -- CP-element group 586: 	575 
    -- CP-element group 586: successors 
    -- CP-element group 586: 	591 
    -- CP-element group 586:  members (3) 
      -- CP-element group 586: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4095_Update/ca
      -- CP-element group 586: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4095_Update/$exit
      -- CP-element group 586: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4095_update_completed_
      -- 
    ca_8882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 586_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4095_inst_ack_1, ack => zeropad3D_CP_2152_elements(586)); -- 
    -- CP-element group 587:  transition  input  bypass 
    -- CP-element group 587: predecessors 
    -- CP-element group 587: 	575 
    -- CP-element group 587: successors 
    -- CP-element group 587:  members (5) 
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_sample_completed_
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Sample/word_access_start/word_0/ra
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Sample/word_access_start/word_0/$exit
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Sample/word_access_start/$exit
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Sample/$exit
      -- 
    ra_8899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 587_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4098_load_0_ack_0, ack => zeropad3D_CP_2152_elements(587)); -- 
    -- CP-element group 588:  transition  input  output  bypass 
    -- CP-element group 588: predecessors 
    -- CP-element group 588: 	575 
    -- CP-element group 588: successors 
    -- CP-element group 588: 	589 
    -- CP-element group 588:  members (12) 
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_update_completed_
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4102_Sample/rr
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4102_Sample/$entry
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4102_sample_start_
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Update/LOAD_row_high_4098_Merge/merge_ack
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Update/LOAD_row_high_4098_Merge/merge_req
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Update/LOAD_row_high_4098_Merge/$exit
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Update/LOAD_row_high_4098_Merge/$entry
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Update/word_access_complete/word_0/ca
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Update/word_access_complete/word_0/$exit
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Update/word_access_complete/$exit
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/LOAD_row_high_4098_Update/$exit
      -- 
    ca_8910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 588_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4098_load_0_ack_1, ack => zeropad3D_CP_2152_elements(588)); -- 
    rr_8923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(588), ack => type_cast_4102_inst_req_0); -- 
    -- CP-element group 589:  transition  input  bypass 
    -- CP-element group 589: predecessors 
    -- CP-element group 589: 	588 
    -- CP-element group 589: successors 
    -- CP-element group 589:  members (3) 
      -- CP-element group 589: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4102_Sample/ra
      -- CP-element group 589: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4102_Sample/$exit
      -- CP-element group 589: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4102_sample_completed_
      -- 
    ra_8924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 589_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4102_inst_ack_0, ack => zeropad3D_CP_2152_elements(589)); -- 
    -- CP-element group 590:  transition  input  bypass 
    -- CP-element group 590: predecessors 
    -- CP-element group 590: 	575 
    -- CP-element group 590: successors 
    -- CP-element group 590: 	591 
    -- CP-element group 590:  members (3) 
      -- CP-element group 590: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4102_Update/ca
      -- CP-element group 590: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4102_Update/$exit
      -- CP-element group 590: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/type_cast_4102_update_completed_
      -- 
    ca_8929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 590_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4102_inst_ack_1, ack => zeropad3D_CP_2152_elements(590)); -- 
    -- CP-element group 591:  branch  join  transition  place  output  bypass 
    -- CP-element group 591: predecessors 
    -- CP-element group 591: 	586 
    -- CP-element group 591: 	590 
    -- CP-element group 591: successors 
    -- CP-element group 591: 	592 
    -- CP-element group 591: 	593 
    -- CP-element group 591:  members (10) 
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125__exit__
      -- CP-element group 591: 	 branch_block_stmt_714/if_stmt_4126__entry__
      -- CP-element group 591: 	 branch_block_stmt_714/if_stmt_4126_eval_test/$entry
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_4054_to_assign_stmt_4125/$exit
      -- CP-element group 591: 	 branch_block_stmt_714/if_stmt_4126_eval_test/$exit
      -- CP-element group 591: 	 branch_block_stmt_714/if_stmt_4126_eval_test/branch_req
      -- CP-element group 591: 	 branch_block_stmt_714/if_stmt_4126_if_link/$entry
      -- CP-element group 591: 	 branch_block_stmt_714/if_stmt_4126_dead_link/$entry
      -- CP-element group 591: 	 branch_block_stmt_714/R_cmp1270_4127_place
      -- CP-element group 591: 	 branch_block_stmt_714/if_stmt_4126_else_link/$entry
      -- 
    branch_req_8937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(591), ack => if_stmt_4126_branch_req_0); -- 
    zeropad3D_cp_element_group_591: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_591"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(586) & zeropad3D_CP_2152_elements(590);
      gj_zeropad3D_cp_element_group_591 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(591), clk => clk, reset => reset); --
    end block;
    -- CP-element group 592:  fork  transition  place  input  output  bypass 
    -- CP-element group 592: predecessors 
    -- CP-element group 592: 	591 
    -- CP-element group 592: successors 
    -- CP-element group 592: 	1116 
    -- CP-element group 592: 	1117 
    -- CP-element group 592: 	1119 
    -- CP-element group 592: 	1120 
    -- CP-element group 592:  members (20) 
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280
      -- CP-element group 592: 	 branch_block_stmt_714/if_stmt_4126_if_link/$exit
      -- CP-element group 592: 	 branch_block_stmt_714/if_stmt_4126_if_link/if_choice_transition
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/$entry
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/$entry
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/$entry
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/type_cast_4158/$entry
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/type_cast_4158/SplitProtocol/$entry
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/type_cast_4158/SplitProtocol/Sample/$entry
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/type_cast_4158/SplitProtocol/Sample/rr
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/type_cast_4158/SplitProtocol/Update/$entry
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/type_cast_4158/SplitProtocol/Update/cr
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/$entry
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/$entry
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/type_cast_4162/$entry
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/type_cast_4162/SplitProtocol/$entry
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/type_cast_4162/SplitProtocol/Sample/$entry
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/type_cast_4162/SplitProtocol/Sample/rr
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/type_cast_4162/SplitProtocol/Update/$entry
      -- CP-element group 592: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/type_cast_4162/SplitProtocol/Update/cr
      -- 
    if_choice_transition_8942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 592_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4126_branch_ack_1, ack => zeropad3D_CP_2152_elements(592)); -- 
    rr_13470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(592), ack => type_cast_4158_inst_req_0); -- 
    cr_13475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(592), ack => type_cast_4158_inst_req_1); -- 
    rr_13493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(592), ack => type_cast_4162_inst_req_0); -- 
    cr_13498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(592), ack => type_cast_4162_inst_req_1); -- 
    -- CP-element group 593:  fork  transition  place  input  output  bypass 
    -- CP-element group 593: predecessors 
    -- CP-element group 593: 	591 
    -- CP-element group 593: successors 
    -- CP-element group 593: 	1093 
    -- CP-element group 593: 	1094 
    -- CP-element group 593: 	1095 
    -- CP-element group 593: 	1097 
    -- CP-element group 593: 	1098 
    -- CP-element group 593:  members (22) 
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279
      -- CP-element group 593: 	 branch_block_stmt_714/if_stmt_4126_else_link/else_choice_transition
      -- CP-element group 593: 	 branch_block_stmt_714/if_stmt_4126_else_link/$exit
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4133/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4145/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4145/SplitProtocol/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4145/SplitProtocol/Sample/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4145/SplitProtocol/Sample/rr
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4145/SplitProtocol/Update/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4145/SplitProtocol/Update/cr
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4151/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4151/SplitProtocol/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4151/SplitProtocol/Sample/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4151/SplitProtocol/Sample/rr
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4151/SplitProtocol/Update/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4151/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 593_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4126_branch_ack_0, ack => zeropad3D_CP_2152_elements(593)); -- 
    rr_13342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(593), ack => type_cast_4145_inst_req_0); -- 
    cr_13347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(593), ack => type_cast_4145_inst_req_1); -- 
    rr_13365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(593), ack => type_cast_4151_inst_req_0); -- 
    cr_13370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(593), ack => type_cast_4151_inst_req_1); -- 
    -- CP-element group 594:  transition  input  bypass 
    -- CP-element group 594: predecessors 
    -- CP-element group 594: 	1125 
    -- CP-element group 594: successors 
    -- CP-element group 594:  members (3) 
      -- CP-element group 594: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4166_Sample/ra
      -- CP-element group 594: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4166_Sample/$exit
      -- CP-element group 594: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4166_sample_completed_
      -- 
    ra_8960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 594_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4166_inst_ack_0, ack => zeropad3D_CP_2152_elements(594)); -- 
    -- CP-element group 595:  transition  input  bypass 
    -- CP-element group 595: predecessors 
    -- CP-element group 595: 	1125 
    -- CP-element group 595: successors 
    -- CP-element group 595: 	608 
    -- CP-element group 595:  members (3) 
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4166_Update/ca
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4166_Update/$exit
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4166_update_completed_
      -- 
    ca_8965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 595_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4166_inst_ack_1, ack => zeropad3D_CP_2152_elements(595)); -- 
    -- CP-element group 596:  transition  input  bypass 
    -- CP-element group 596: predecessors 
    -- CP-element group 596: 	1125 
    -- CP-element group 596: successors 
    -- CP-element group 596:  members (5) 
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Sample/word_access_start/$exit
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Sample/word_access_start/word_0/$exit
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Sample/$exit
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Sample/word_access_start/word_0/ra
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_sample_completed_
      -- 
    ra_8982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 596_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_4181_load_0_ack_0, ack => zeropad3D_CP_2152_elements(596)); -- 
    -- CP-element group 597:  transition  input  output  bypass 
    -- CP-element group 597: predecessors 
    -- CP-element group 597: 	1125 
    -- CP-element group 597: successors 
    -- CP-element group 597: 	606 
    -- CP-element group 597:  members (12) 
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Update/$exit
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Update/word_access_complete/word_0/ca
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Update/word_access_complete/$exit
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Update/word_access_complete/word_0/$exit
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_update_completed_
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Update/LOAD_pad_4181_Merge/$entry
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Update/LOAD_pad_4181_Merge/merge_ack
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Update/LOAD_pad_4181_Merge/merge_req
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Update/LOAD_pad_4181_Merge/$exit
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4251_sample_start_
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4251_Sample/$entry
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4251_Sample/rr
      -- 
    ca_8993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 597_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_4181_load_0_ack_1, ack => zeropad3D_CP_2152_elements(597)); -- 
    rr_9153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(597), ack => type_cast_4251_inst_req_0); -- 
    -- CP-element group 598:  transition  input  bypass 
    -- CP-element group 598: predecessors 
    -- CP-element group 598: 	1125 
    -- CP-element group 598: successors 
    -- CP-element group 598:  members (5) 
      -- CP-element group 598: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Sample/word_access_start/word_0/ra
      -- CP-element group 598: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Sample/word_access_start/word_0/$exit
      -- CP-element group 598: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Sample/word_access_start/$exit
      -- CP-element group 598: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Sample/$exit
      -- CP-element group 598: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_sample_completed_
      -- 
    ra_9015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 598_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_4184_load_0_ack_0, ack => zeropad3D_CP_2152_elements(598)); -- 
    -- CP-element group 599:  transition  input  output  bypass 
    -- CP-element group 599: predecessors 
    -- CP-element group 599: 	1125 
    -- CP-element group 599: successors 
    -- CP-element group 599: 	604 
    -- CP-element group 599:  members (12) 
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Update/LOAD_depth_high_4184_Merge/merge_ack
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Update/LOAD_depth_high_4184_Merge/merge_req
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Update/LOAD_depth_high_4184_Merge/$exit
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Update/LOAD_depth_high_4184_Merge/$entry
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Update/word_access_complete/word_0/ca
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Update/word_access_complete/word_0/$exit
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Update/word_access_complete/$exit
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Update/$exit
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_update_completed_
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4212_sample_start_
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4212_Sample/$entry
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4212_Sample/rr
      -- 
    ca_9026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 599_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_4184_load_0_ack_1, ack => zeropad3D_CP_2152_elements(599)); -- 
    rr_9139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(599), ack => type_cast_4212_inst_req_0); -- 
    -- CP-element group 600:  transition  input  bypass 
    -- CP-element group 600: predecessors 
    -- CP-element group 600: 	1125 
    -- CP-element group 600: successors 
    -- CP-element group 600:  members (5) 
      -- CP-element group 600: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_sample_completed_
      -- CP-element group 600: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Sample/word_access_start/word_0/ra
      -- CP-element group 600: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Sample/word_access_start/word_0/$exit
      -- CP-element group 600: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Sample/word_access_start/$exit
      -- CP-element group 600: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Sample/$exit
      -- 
    ra_9065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 600_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4196_load_0_ack_0, ack => zeropad3D_CP_2152_elements(600)); -- 
    -- CP-element group 601:  transition  input  bypass 
    -- CP-element group 601: predecessors 
    -- CP-element group 601: 	1125 
    -- CP-element group 601: successors 
    -- CP-element group 601: 	608 
    -- CP-element group 601:  members (9) 
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_update_completed_
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Update/word_access_complete/word_0/$exit
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Update/word_access_complete/$exit
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Update/$exit
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Update/word_access_complete/word_0/ca
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Update/ptr_deref_4196_Merge/$entry
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Update/ptr_deref_4196_Merge/$exit
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Update/ptr_deref_4196_Merge/merge_req
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Update/ptr_deref_4196_Merge/merge_ack
      -- 
    ca_9076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 601_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4196_load_0_ack_1, ack => zeropad3D_CP_2152_elements(601)); -- 
    -- CP-element group 602:  transition  input  bypass 
    -- CP-element group 602: predecessors 
    -- CP-element group 602: 	1125 
    -- CP-element group 602: successors 
    -- CP-element group 602:  members (5) 
      -- CP-element group 602: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_sample_completed_
      -- CP-element group 602: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Sample/$exit
      -- CP-element group 602: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Sample/word_access_start/$exit
      -- CP-element group 602: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Sample/word_access_start/word_0/$exit
      -- CP-element group 602: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Sample/word_access_start/word_0/ra
      -- 
    ra_9115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 602_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4208_load_0_ack_0, ack => zeropad3D_CP_2152_elements(602)); -- 
    -- CP-element group 603:  transition  input  bypass 
    -- CP-element group 603: predecessors 
    -- CP-element group 603: 	1125 
    -- CP-element group 603: successors 
    -- CP-element group 603: 	608 
    -- CP-element group 603:  members (9) 
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_update_completed_
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Update/$exit
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Update/word_access_complete/$exit
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Update/word_access_complete/word_0/$exit
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Update/word_access_complete/word_0/ca
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Update/ptr_deref_4208_Merge/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Update/ptr_deref_4208_Merge/$exit
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Update/ptr_deref_4208_Merge/merge_req
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Update/ptr_deref_4208_Merge/merge_ack
      -- 
    ca_9126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 603_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4208_load_0_ack_1, ack => zeropad3D_CP_2152_elements(603)); -- 
    -- CP-element group 604:  transition  input  bypass 
    -- CP-element group 604: predecessors 
    -- CP-element group 604: 	599 
    -- CP-element group 604: successors 
    -- CP-element group 604:  members (3) 
      -- CP-element group 604: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4212_sample_completed_
      -- CP-element group 604: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4212_Sample/$exit
      -- CP-element group 604: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4212_Sample/ra
      -- 
    ra_9140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 604_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4212_inst_ack_0, ack => zeropad3D_CP_2152_elements(604)); -- 
    -- CP-element group 605:  transition  input  bypass 
    -- CP-element group 605: predecessors 
    -- CP-element group 605: 	1125 
    -- CP-element group 605: successors 
    -- CP-element group 605: 	608 
    -- CP-element group 605:  members (3) 
      -- CP-element group 605: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4212_update_completed_
      -- CP-element group 605: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4212_Update/$exit
      -- CP-element group 605: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4212_Update/ca
      -- 
    ca_9145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 605_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4212_inst_ack_1, ack => zeropad3D_CP_2152_elements(605)); -- 
    -- CP-element group 606:  transition  input  bypass 
    -- CP-element group 606: predecessors 
    -- CP-element group 606: 	597 
    -- CP-element group 606: successors 
    -- CP-element group 606:  members (3) 
      -- CP-element group 606: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4251_sample_completed_
      -- CP-element group 606: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4251_Sample/$exit
      -- CP-element group 606: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4251_Sample/ra
      -- 
    ra_9154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 606_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4251_inst_ack_0, ack => zeropad3D_CP_2152_elements(606)); -- 
    -- CP-element group 607:  transition  input  bypass 
    -- CP-element group 607: predecessors 
    -- CP-element group 607: 	1125 
    -- CP-element group 607: successors 
    -- CP-element group 607: 	608 
    -- CP-element group 607:  members (3) 
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4251_update_completed_
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4251_Update/$exit
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4251_Update/ca
      -- 
    ca_9159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 607_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4251_inst_ack_1, ack => zeropad3D_CP_2152_elements(607)); -- 
    -- CP-element group 608:  join  fork  transition  place  output  bypass 
    -- CP-element group 608: predecessors 
    -- CP-element group 608: 	595 
    -- CP-element group 608: 	601 
    -- CP-element group 608: 	603 
    -- CP-element group 608: 	605 
    -- CP-element group 608: 	607 
    -- CP-element group 608: successors 
    -- CP-element group 608: 	1136 
    -- CP-element group 608: 	1137 
    -- CP-element group 608: 	1138 
    -- CP-element group 608: 	1140 
    -- CP-element group 608:  members (16) 
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341
      -- CP-element group 608: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293__exit__
      -- CP-element group 608: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/$exit
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/$entry
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4296/$entry
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/$entry
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/$entry
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/$entry
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4306/$entry
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4306/SplitProtocol/$entry
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4306/SplitProtocol/Sample/$entry
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4306/SplitProtocol/Sample/rr
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4306/SplitProtocol/Update/$entry
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4306/SplitProtocol/Update/cr
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4309/$entry
      -- CP-element group 608: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/$entry
      -- 
    rr_13605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(608), ack => type_cast_4306_inst_req_0); -- 
    cr_13610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(608), ack => type_cast_4306_inst_req_1); -- 
    zeropad3D_cp_element_group_608: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_608"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(595) & zeropad3D_CP_2152_elements(601) & zeropad3D_CP_2152_elements(603) & zeropad3D_CP_2152_elements(605) & zeropad3D_CP_2152_elements(607);
      gj_zeropad3D_cp_element_group_608 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(608), clk => clk, reset => reset); --
    end block;
    -- CP-element group 609:  transition  input  bypass 
    -- CP-element group 609: predecessors 
    -- CP-element group 609: 	1146 
    -- CP-element group 609: successors 
    -- CP-element group 609:  members (3) 
      -- CP-element group 609: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/type_cast_4320_sample_completed_
      -- CP-element group 609: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/type_cast_4320_Sample/$exit
      -- CP-element group 609: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/type_cast_4320_Sample/ra
      -- 
    ra_9171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 609_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4320_inst_ack_0, ack => zeropad3D_CP_2152_elements(609)); -- 
    -- CP-element group 610:  branch  transition  place  input  output  bypass 
    -- CP-element group 610: predecessors 
    -- CP-element group 610: 	1146 
    -- CP-element group 610: successors 
    -- CP-element group 610: 	611 
    -- CP-element group 610: 	612 
    -- CP-element group 610:  members (13) 
      -- CP-element group 610: 	 branch_block_stmt_714/if_stmt_4329__entry__
      -- CP-element group 610: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328__exit__
      -- CP-element group 610: 	 branch_block_stmt_714/R_cmp1346_4330_place
      -- CP-element group 610: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/$exit
      -- CP-element group 610: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/type_cast_4320_update_completed_
      -- CP-element group 610: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/type_cast_4320_Update/$exit
      -- CP-element group 610: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/type_cast_4320_Update/ca
      -- CP-element group 610: 	 branch_block_stmt_714/if_stmt_4329_dead_link/$entry
      -- CP-element group 610: 	 branch_block_stmt_714/if_stmt_4329_eval_test/$entry
      -- CP-element group 610: 	 branch_block_stmt_714/if_stmt_4329_eval_test/$exit
      -- CP-element group 610: 	 branch_block_stmt_714/if_stmt_4329_eval_test/branch_req
      -- CP-element group 610: 	 branch_block_stmt_714/if_stmt_4329_if_link/$entry
      -- CP-element group 610: 	 branch_block_stmt_714/if_stmt_4329_else_link/$entry
      -- 
    ca_9176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 610_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4320_inst_ack_1, ack => zeropad3D_CP_2152_elements(610)); -- 
    branch_req_9184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(610), ack => if_stmt_4329_branch_req_0); -- 
    -- CP-element group 611:  transition  place  input  bypass 
    -- CP-element group 611: predecessors 
    -- CP-element group 611: 	610 
    -- CP-element group 611: successors 
    -- CP-element group 611: 	1147 
    -- CP-element group 611:  members (5) 
      -- CP-element group 611: 	 branch_block_stmt_714/whilex_xbody1341_ifx_xthen1376
      -- CP-element group 611: 	 branch_block_stmt_714/if_stmt_4329_if_link/$exit
      -- CP-element group 611: 	 branch_block_stmt_714/if_stmt_4329_if_link/if_choice_transition
      -- CP-element group 611: 	 branch_block_stmt_714/whilex_xbody1341_ifx_xthen1376_PhiReq/$entry
      -- CP-element group 611: 	 branch_block_stmt_714/whilex_xbody1341_ifx_xthen1376_PhiReq/$exit
      -- 
    if_choice_transition_9189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 611_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4329_branch_ack_1, ack => zeropad3D_CP_2152_elements(611)); -- 
    -- CP-element group 612:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 612: predecessors 
    -- CP-element group 612: 	610 
    -- CP-element group 612: successors 
    -- CP-element group 612: 	613 
    -- CP-element group 612: 	614 
    -- CP-element group 612: 	616 
    -- CP-element group 612:  members (27) 
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354__entry__
      -- CP-element group 612: 	 branch_block_stmt_714/merge_stmt_4335__exit__
      -- CP-element group 612: 	 branch_block_stmt_714/whilex_xbody1341_lorx_xlhsx_xfalse1348
      -- CP-element group 612: 	 branch_block_stmt_714/if_stmt_4329_else_link/$exit
      -- CP-element group 612: 	 branch_block_stmt_714/if_stmt_4329_else_link/else_choice_transition
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/$entry
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_sample_start_
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_update_start_
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_word_address_calculated
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_root_address_calculated
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Sample/$entry
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Sample/word_access_start/$entry
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Sample/word_access_start/word_0/$entry
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Sample/word_access_start/word_0/rr
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Update/$entry
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Update/word_access_complete/$entry
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Update/word_access_complete/word_0/$entry
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Update/word_access_complete/word_0/cr
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/type_cast_4341_update_start_
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/type_cast_4341_Update/$entry
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/type_cast_4341_Update/cr
      -- CP-element group 612: 	 branch_block_stmt_714/whilex_xbody1341_lorx_xlhsx_xfalse1348_PhiReq/$entry
      -- CP-element group 612: 	 branch_block_stmt_714/whilex_xbody1341_lorx_xlhsx_xfalse1348_PhiReq/$exit
      -- CP-element group 612: 	 branch_block_stmt_714/merge_stmt_4335_PhiReqMerge
      -- CP-element group 612: 	 branch_block_stmt_714/merge_stmt_4335_PhiAck/$entry
      -- CP-element group 612: 	 branch_block_stmt_714/merge_stmt_4335_PhiAck/$exit
      -- CP-element group 612: 	 branch_block_stmt_714/merge_stmt_4335_PhiAck/dummy
      -- 
    else_choice_transition_9193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 612_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4329_branch_ack_0, ack => zeropad3D_CP_2152_elements(612)); -- 
    rr_9214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(612), ack => LOAD_row_high_4337_load_0_req_0); -- 
    cr_9225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(612), ack => LOAD_row_high_4337_load_0_req_1); -- 
    cr_9244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(612), ack => type_cast_4341_inst_req_1); -- 
    -- CP-element group 613:  transition  input  bypass 
    -- CP-element group 613: predecessors 
    -- CP-element group 613: 	612 
    -- CP-element group 613: successors 
    -- CP-element group 613:  members (5) 
      -- CP-element group 613: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_sample_completed_
      -- CP-element group 613: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Sample/$exit
      -- CP-element group 613: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Sample/word_access_start/$exit
      -- CP-element group 613: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Sample/word_access_start/word_0/$exit
      -- CP-element group 613: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Sample/word_access_start/word_0/ra
      -- 
    ra_9215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 613_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4337_load_0_ack_0, ack => zeropad3D_CP_2152_elements(613)); -- 
    -- CP-element group 614:  transition  input  output  bypass 
    -- CP-element group 614: predecessors 
    -- CP-element group 614: 	612 
    -- CP-element group 614: successors 
    -- CP-element group 614: 	615 
    -- CP-element group 614:  members (12) 
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_update_completed_
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Update/$exit
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Update/word_access_complete/$exit
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Update/word_access_complete/word_0/$exit
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Update/word_access_complete/word_0/ca
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Update/LOAD_row_high_4337_Merge/$entry
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Update/LOAD_row_high_4337_Merge/$exit
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Update/LOAD_row_high_4337_Merge/merge_req
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/LOAD_row_high_4337_Update/LOAD_row_high_4337_Merge/merge_ack
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/type_cast_4341_sample_start_
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/type_cast_4341_Sample/$entry
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/type_cast_4341_Sample/rr
      -- 
    ca_9226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 614_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4337_load_0_ack_1, ack => zeropad3D_CP_2152_elements(614)); -- 
    rr_9239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(614), ack => type_cast_4341_inst_req_0); -- 
    -- CP-element group 615:  transition  input  bypass 
    -- CP-element group 615: predecessors 
    -- CP-element group 615: 	614 
    -- CP-element group 615: successors 
    -- CP-element group 615:  members (3) 
      -- CP-element group 615: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/type_cast_4341_sample_completed_
      -- CP-element group 615: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/type_cast_4341_Sample/$exit
      -- CP-element group 615: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/type_cast_4341_Sample/ra
      -- 
    ra_9240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 615_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4341_inst_ack_0, ack => zeropad3D_CP_2152_elements(615)); -- 
    -- CP-element group 616:  branch  transition  place  input  output  bypass 
    -- CP-element group 616: predecessors 
    -- CP-element group 616: 	612 
    -- CP-element group 616: successors 
    -- CP-element group 616: 	617 
    -- CP-element group 616: 	618 
    -- CP-element group 616:  members (13) 
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354__exit__
      -- CP-element group 616: 	 branch_block_stmt_714/if_stmt_4355__entry__
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/$exit
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/type_cast_4341_update_completed_
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/type_cast_4341_Update/$exit
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4338_to_assign_stmt_4354/type_cast_4341_Update/ca
      -- CP-element group 616: 	 branch_block_stmt_714/if_stmt_4355_dead_link/$entry
      -- CP-element group 616: 	 branch_block_stmt_714/if_stmt_4355_eval_test/$entry
      -- CP-element group 616: 	 branch_block_stmt_714/if_stmt_4355_eval_test/$exit
      -- CP-element group 616: 	 branch_block_stmt_714/if_stmt_4355_eval_test/branch_req
      -- CP-element group 616: 	 branch_block_stmt_714/R_cmp1356_4356_place
      -- CP-element group 616: 	 branch_block_stmt_714/if_stmt_4355_if_link/$entry
      -- CP-element group 616: 	 branch_block_stmt_714/if_stmt_4355_else_link/$entry
      -- 
    ca_9245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 616_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4341_inst_ack_1, ack => zeropad3D_CP_2152_elements(616)); -- 
    branch_req_9253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(616), ack => if_stmt_4355_branch_req_0); -- 
    -- CP-element group 617:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 617: predecessors 
    -- CP-element group 617: 	616 
    -- CP-element group 617: successors 
    -- CP-element group 617: 	619 
    -- CP-element group 617: 	620 
    -- CP-element group 617:  members (18) 
      -- CP-element group 617: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373__entry__
      -- CP-element group 617: 	 branch_block_stmt_714/merge_stmt_4361__exit__
      -- CP-element group 617: 	 branch_block_stmt_714/if_stmt_4355_if_link/$exit
      -- CP-element group 617: 	 branch_block_stmt_714/if_stmt_4355_if_link/if_choice_transition
      -- CP-element group 617: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1348_lorx_xlhsx_xfalse1358
      -- CP-element group 617: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/$entry
      -- CP-element group 617: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/type_cast_4365_sample_start_
      -- CP-element group 617: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/type_cast_4365_update_start_
      -- CP-element group 617: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/type_cast_4365_Sample/$entry
      -- CP-element group 617: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/type_cast_4365_Sample/rr
      -- CP-element group 617: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/type_cast_4365_Update/$entry
      -- CP-element group 617: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/type_cast_4365_Update/cr
      -- CP-element group 617: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1348_lorx_xlhsx_xfalse1358_PhiReq/$entry
      -- CP-element group 617: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1348_lorx_xlhsx_xfalse1358_PhiReq/$exit
      -- CP-element group 617: 	 branch_block_stmt_714/merge_stmt_4361_PhiReqMerge
      -- CP-element group 617: 	 branch_block_stmt_714/merge_stmt_4361_PhiAck/$entry
      -- CP-element group 617: 	 branch_block_stmt_714/merge_stmt_4361_PhiAck/$exit
      -- CP-element group 617: 	 branch_block_stmt_714/merge_stmt_4361_PhiAck/dummy
      -- 
    if_choice_transition_9258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 617_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4355_branch_ack_1, ack => zeropad3D_CP_2152_elements(617)); -- 
    rr_9275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(617), ack => type_cast_4365_inst_req_0); -- 
    cr_9280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(617), ack => type_cast_4365_inst_req_1); -- 
    -- CP-element group 618:  transition  place  input  bypass 
    -- CP-element group 618: predecessors 
    -- CP-element group 618: 	616 
    -- CP-element group 618: successors 
    -- CP-element group 618: 	1147 
    -- CP-element group 618:  members (5) 
      -- CP-element group 618: 	 branch_block_stmt_714/if_stmt_4355_else_link/$exit
      -- CP-element group 618: 	 branch_block_stmt_714/if_stmt_4355_else_link/else_choice_transition
      -- CP-element group 618: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1348_ifx_xthen1376
      -- CP-element group 618: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1348_ifx_xthen1376_PhiReq/$entry
      -- CP-element group 618: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1348_ifx_xthen1376_PhiReq/$exit
      -- 
    else_choice_transition_9262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 618_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4355_branch_ack_0, ack => zeropad3D_CP_2152_elements(618)); -- 
    -- CP-element group 619:  transition  input  bypass 
    -- CP-element group 619: predecessors 
    -- CP-element group 619: 	617 
    -- CP-element group 619: successors 
    -- CP-element group 619:  members (3) 
      -- CP-element group 619: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/type_cast_4365_sample_completed_
      -- CP-element group 619: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/type_cast_4365_Sample/$exit
      -- CP-element group 619: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/type_cast_4365_Sample/ra
      -- 
    ra_9276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 619_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4365_inst_ack_0, ack => zeropad3D_CP_2152_elements(619)); -- 
    -- CP-element group 620:  branch  transition  place  input  output  bypass 
    -- CP-element group 620: predecessors 
    -- CP-element group 620: 	617 
    -- CP-element group 620: successors 
    -- CP-element group 620: 	621 
    -- CP-element group 620: 	622 
    -- CP-element group 620:  members (13) 
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373__exit__
      -- CP-element group 620: 	 branch_block_stmt_714/if_stmt_4374__entry__
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/$exit
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/type_cast_4365_update_completed_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/type_cast_4365_Update/$exit
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4366_to_assign_stmt_4373/type_cast_4365_Update/ca
      -- CP-element group 620: 	 branch_block_stmt_714/if_stmt_4374_dead_link/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/if_stmt_4374_eval_test/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/if_stmt_4374_eval_test/$exit
      -- CP-element group 620: 	 branch_block_stmt_714/if_stmt_4374_eval_test/branch_req
      -- CP-element group 620: 	 branch_block_stmt_714/R_cmp1363_4375_place
      -- CP-element group 620: 	 branch_block_stmt_714/if_stmt_4374_if_link/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/if_stmt_4374_else_link/$entry
      -- 
    ca_9281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 620_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4365_inst_ack_1, ack => zeropad3D_CP_2152_elements(620)); -- 
    branch_req_9289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => if_stmt_4374_branch_req_0); -- 
    -- CP-element group 621:  transition  place  input  bypass 
    -- CP-element group 621: predecessors 
    -- CP-element group 621: 	620 
    -- CP-element group 621: successors 
    -- CP-element group 621: 	1147 
    -- CP-element group 621:  members (5) 
      -- CP-element group 621: 	 branch_block_stmt_714/if_stmt_4374_if_link/$exit
      -- CP-element group 621: 	 branch_block_stmt_714/if_stmt_4374_if_link/if_choice_transition
      -- CP-element group 621: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1358_ifx_xthen1376
      -- CP-element group 621: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1358_ifx_xthen1376_PhiReq/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1358_ifx_xthen1376_PhiReq/$exit
      -- 
    if_choice_transition_9294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 621_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4374_branch_ack_1, ack => zeropad3D_CP_2152_elements(621)); -- 
    -- CP-element group 622:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 622: predecessors 
    -- CP-element group 622: 	620 
    -- CP-element group 622: successors 
    -- CP-element group 622: 	623 
    -- CP-element group 622: 	624 
    -- CP-element group 622: 	626 
    -- CP-element group 622:  members (27) 
      -- CP-element group 622: 	 branch_block_stmt_714/merge_stmt_4380__exit__
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405__entry__
      -- CP-element group 622: 	 branch_block_stmt_714/if_stmt_4374_else_link/$exit
      -- CP-element group 622: 	 branch_block_stmt_714/if_stmt_4374_else_link/else_choice_transition
      -- CP-element group 622: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1358_lorx_xlhsx_xfalse1365
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/$entry
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_sample_start_
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_update_start_
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_word_address_calculated
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_root_address_calculated
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Sample/$entry
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Sample/word_access_start/$entry
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Sample/word_access_start/word_0/$entry
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Sample/word_access_start/word_0/rr
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Update/$entry
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Update/word_access_complete/$entry
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Update/word_access_complete/word_0/$entry
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Update/word_access_complete/word_0/cr
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/type_cast_4386_update_start_
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/type_cast_4386_Update/$entry
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/type_cast_4386_Update/cr
      -- CP-element group 622: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1358_lorx_xlhsx_xfalse1365_PhiReq/$entry
      -- CP-element group 622: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1358_lorx_xlhsx_xfalse1365_PhiReq/$exit
      -- CP-element group 622: 	 branch_block_stmt_714/merge_stmt_4380_PhiReqMerge
      -- CP-element group 622: 	 branch_block_stmt_714/merge_stmt_4380_PhiAck/$entry
      -- CP-element group 622: 	 branch_block_stmt_714/merge_stmt_4380_PhiAck/$exit
      -- CP-element group 622: 	 branch_block_stmt_714/merge_stmt_4380_PhiAck/dummy
      -- 
    else_choice_transition_9298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 622_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4374_branch_ack_0, ack => zeropad3D_CP_2152_elements(622)); -- 
    rr_9319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(622), ack => LOAD_col_high_4382_load_0_req_0); -- 
    cr_9330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(622), ack => LOAD_col_high_4382_load_0_req_1); -- 
    cr_9349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(622), ack => type_cast_4386_inst_req_1); -- 
    -- CP-element group 623:  transition  input  bypass 
    -- CP-element group 623: predecessors 
    -- CP-element group 623: 	622 
    -- CP-element group 623: successors 
    -- CP-element group 623:  members (5) 
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_sample_completed_
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Sample/$exit
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Sample/word_access_start/$exit
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Sample/word_access_start/word_0/$exit
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Sample/word_access_start/word_0/ra
      -- 
    ra_9320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 623_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4382_load_0_ack_0, ack => zeropad3D_CP_2152_elements(623)); -- 
    -- CP-element group 624:  transition  input  output  bypass 
    -- CP-element group 624: predecessors 
    -- CP-element group 624: 	622 
    -- CP-element group 624: successors 
    -- CP-element group 624: 	625 
    -- CP-element group 624:  members (12) 
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_update_completed_
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Update/$exit
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Update/word_access_complete/$exit
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Update/word_access_complete/word_0/$exit
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Update/word_access_complete/word_0/ca
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Update/LOAD_col_high_4382_Merge/$entry
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Update/LOAD_col_high_4382_Merge/$exit
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Update/LOAD_col_high_4382_Merge/merge_req
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/LOAD_col_high_4382_Update/LOAD_col_high_4382_Merge/merge_ack
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/type_cast_4386_sample_start_
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/type_cast_4386_Sample/$entry
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/type_cast_4386_Sample/rr
      -- 
    ca_9331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 624_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4382_load_0_ack_1, ack => zeropad3D_CP_2152_elements(624)); -- 
    rr_9344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(624), ack => type_cast_4386_inst_req_0); -- 
    -- CP-element group 625:  transition  input  bypass 
    -- CP-element group 625: predecessors 
    -- CP-element group 625: 	624 
    -- CP-element group 625: successors 
    -- CP-element group 625:  members (3) 
      -- CP-element group 625: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/type_cast_4386_sample_completed_
      -- CP-element group 625: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/type_cast_4386_Sample/$exit
      -- CP-element group 625: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/type_cast_4386_Sample/ra
      -- 
    ra_9345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 625_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4386_inst_ack_0, ack => zeropad3D_CP_2152_elements(625)); -- 
    -- CP-element group 626:  branch  transition  place  input  output  bypass 
    -- CP-element group 626: predecessors 
    -- CP-element group 626: 	622 
    -- CP-element group 626: successors 
    -- CP-element group 626: 	627 
    -- CP-element group 626: 	628 
    -- CP-element group 626:  members (13) 
      -- CP-element group 626: 	 branch_block_stmt_714/if_stmt_4406__entry__
      -- CP-element group 626: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405__exit__
      -- CP-element group 626: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/$exit
      -- CP-element group 626: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/type_cast_4386_update_completed_
      -- CP-element group 626: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/type_cast_4386_Update/$exit
      -- CP-element group 626: 	 branch_block_stmt_714/assign_stmt_4383_to_assign_stmt_4405/type_cast_4386_Update/ca
      -- CP-element group 626: 	 branch_block_stmt_714/if_stmt_4406_dead_link/$entry
      -- CP-element group 626: 	 branch_block_stmt_714/if_stmt_4406_eval_test/$entry
      -- CP-element group 626: 	 branch_block_stmt_714/if_stmt_4406_eval_test/$exit
      -- CP-element group 626: 	 branch_block_stmt_714/if_stmt_4406_eval_test/branch_req
      -- CP-element group 626: 	 branch_block_stmt_714/R_cmp1374_4407_place
      -- CP-element group 626: 	 branch_block_stmt_714/if_stmt_4406_if_link/$entry
      -- CP-element group 626: 	 branch_block_stmt_714/if_stmt_4406_else_link/$entry
      -- 
    ca_9350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 626_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4386_inst_ack_1, ack => zeropad3D_CP_2152_elements(626)); -- 
    branch_req_9358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(626), ack => if_stmt_4406_branch_req_0); -- 
    -- CP-element group 627:  fork  transition  place  input  output  bypass 
    -- CP-element group 627: predecessors 
    -- CP-element group 627: 	626 
    -- CP-element group 627: successors 
    -- CP-element group 627: 	643 
    -- CP-element group 627: 	644 
    -- CP-element group 627: 	646 
    -- CP-element group 627: 	648 
    -- CP-element group 627: 	650 
    -- CP-element group 627: 	652 
    -- CP-element group 627: 	654 
    -- CP-element group 627: 	656 
    -- CP-element group 627: 	658 
    -- CP-element group 627: 	661 
    -- CP-element group 627:  members (46) 
      -- CP-element group 627: 	 branch_block_stmt_714/merge_stmt_4470__exit__
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575__entry__
      -- CP-element group 627: 	 branch_block_stmt_714/if_stmt_4406_if_link/$exit
      -- CP-element group 627: 	 branch_block_stmt_714/if_stmt_4406_if_link/if_choice_transition
      -- CP-element group 627: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1365_ifx_xelse1397
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4474_sample_start_
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4474_update_start_
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4474_Sample/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4474_Sample/rr
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4474_Update/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4474_Update/cr
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4538_update_start_
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4538_Update/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4538_Update/cr
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4545_update_start_
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Update/word_access_complete/word_0/cr
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_final_index_sum_regn_update_start
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_final_index_sum_regn_Update/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_final_index_sum_regn_Update/req
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4545_complete/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4545_complete/req
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_update_start_
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Update/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Update/word_access_complete/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Update/word_access_complete/word_0/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Update/word_access_complete/word_0/cr
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4563_update_start_
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4563_Update/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4563_Update/cr
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4570_update_start_
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Update/word_access_complete/word_0/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_final_index_sum_regn_update_start
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_final_index_sum_regn_Update/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_final_index_sum_regn_Update/req
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Update/word_access_complete/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4570_complete/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4570_complete/req
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_update_start_
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Update/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1365_ifx_xelse1397_PhiReq/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1365_ifx_xelse1397_PhiReq/$exit
      -- CP-element group 627: 	 branch_block_stmt_714/merge_stmt_4470_PhiReqMerge
      -- CP-element group 627: 	 branch_block_stmt_714/merge_stmt_4470_PhiAck/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/merge_stmt_4470_PhiAck/$exit
      -- CP-element group 627: 	 branch_block_stmt_714/merge_stmt_4470_PhiAck/dummy
      -- 
    if_choice_transition_9363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 627_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4406_branch_ack_1, ack => zeropad3D_CP_2152_elements(627)); -- 
    rr_9521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(627), ack => type_cast_4474_inst_req_0); -- 
    cr_9526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(627), ack => type_cast_4474_inst_req_1); -- 
    cr_9540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(627), ack => type_cast_4538_inst_req_1); -- 
    cr_9746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(627), ack => ptr_deref_4573_store_0_req_1); -- 
    req_9571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(627), ack => array_obj_ref_4544_index_offset_req_1); -- 
    req_9586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(627), ack => addr_of_4545_final_reg_req_1); -- 
    cr_9631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(627), ack => ptr_deref_4549_load_0_req_1); -- 
    cr_9650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(627), ack => type_cast_4563_inst_req_1); -- 
    req_9681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(627), ack => array_obj_ref_4569_index_offset_req_1); -- 
    req_9696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(627), ack => addr_of_4570_final_reg_req_1); -- 
    -- CP-element group 628:  transition  place  input  bypass 
    -- CP-element group 628: predecessors 
    -- CP-element group 628: 	626 
    -- CP-element group 628: successors 
    -- CP-element group 628: 	1147 
    -- CP-element group 628:  members (5) 
      -- CP-element group 628: 	 branch_block_stmt_714/if_stmt_4406_else_link/$exit
      -- CP-element group 628: 	 branch_block_stmt_714/if_stmt_4406_else_link/else_choice_transition
      -- CP-element group 628: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1365_ifx_xthen1376
      -- CP-element group 628: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1365_ifx_xthen1376_PhiReq/$entry
      -- CP-element group 628: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1365_ifx_xthen1376_PhiReq/$exit
      -- 
    else_choice_transition_9367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 628_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4406_branch_ack_0, ack => zeropad3D_CP_2152_elements(628)); -- 
    -- CP-element group 629:  transition  input  bypass 
    -- CP-element group 629: predecessors 
    -- CP-element group 629: 	1147 
    -- CP-element group 629: successors 
    -- CP-element group 629:  members (3) 
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4416_sample_completed_
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4416_Sample/$exit
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4416_Sample/ra
      -- 
    ra_9381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 629_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4416_inst_ack_0, ack => zeropad3D_CP_2152_elements(629)); -- 
    -- CP-element group 630:  transition  input  bypass 
    -- CP-element group 630: predecessors 
    -- CP-element group 630: 	1147 
    -- CP-element group 630: successors 
    -- CP-element group 630: 	633 
    -- CP-element group 630:  members (3) 
      -- CP-element group 630: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4416_update_completed_
      -- CP-element group 630: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4416_Update/$exit
      -- CP-element group 630: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4416_Update/ca
      -- 
    ca_9386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 630_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4416_inst_ack_1, ack => zeropad3D_CP_2152_elements(630)); -- 
    -- CP-element group 631:  transition  input  bypass 
    -- CP-element group 631: predecessors 
    -- CP-element group 631: 	1147 
    -- CP-element group 631: successors 
    -- CP-element group 631:  members (3) 
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4421_sample_completed_
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4421_Sample/$exit
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4421_Sample/ra
      -- 
    ra_9395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 631_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4421_inst_ack_0, ack => zeropad3D_CP_2152_elements(631)); -- 
    -- CP-element group 632:  transition  input  bypass 
    -- CP-element group 632: predecessors 
    -- CP-element group 632: 	1147 
    -- CP-element group 632: successors 
    -- CP-element group 632: 	633 
    -- CP-element group 632:  members (3) 
      -- CP-element group 632: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4421_update_completed_
      -- CP-element group 632: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4421_Update/$exit
      -- CP-element group 632: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4421_Update/ca
      -- 
    ca_9400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 632_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4421_inst_ack_1, ack => zeropad3D_CP_2152_elements(632)); -- 
    -- CP-element group 633:  join  transition  output  bypass 
    -- CP-element group 633: predecessors 
    -- CP-element group 633: 	630 
    -- CP-element group 633: 	632 
    -- CP-element group 633: successors 
    -- CP-element group 633: 	634 
    -- CP-element group 633:  members (3) 
      -- CP-element group 633: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4455_sample_start_
      -- CP-element group 633: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4455_Sample/$entry
      -- CP-element group 633: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4455_Sample/rr
      -- 
    rr_9408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(633), ack => type_cast_4455_inst_req_0); -- 
    zeropad3D_cp_element_group_633: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_633"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(630) & zeropad3D_CP_2152_elements(632);
      gj_zeropad3D_cp_element_group_633 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(633), clk => clk, reset => reset); --
    end block;
    -- CP-element group 634:  transition  input  bypass 
    -- CP-element group 634: predecessors 
    -- CP-element group 634: 	633 
    -- CP-element group 634: successors 
    -- CP-element group 634:  members (3) 
      -- CP-element group 634: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4455_sample_completed_
      -- CP-element group 634: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4455_Sample/$exit
      -- CP-element group 634: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4455_Sample/ra
      -- 
    ra_9409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 634_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4455_inst_ack_0, ack => zeropad3D_CP_2152_elements(634)); -- 
    -- CP-element group 635:  transition  input  output  bypass 
    -- CP-element group 635: predecessors 
    -- CP-element group 635: 	1147 
    -- CP-element group 635: successors 
    -- CP-element group 635: 	636 
    -- CP-element group 635:  members (16) 
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4455_update_completed_
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4455_Update/$exit
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4455_Update/ca
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_index_resized_1
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_index_scaled_1
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_index_computed_1
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_index_resize_1/$entry
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_index_resize_1/$exit
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_index_resize_1/index_resize_req
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_index_resize_1/index_resize_ack
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_index_scale_1/$entry
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_index_scale_1/$exit
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_index_scale_1/scale_rename_req
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_index_scale_1/scale_rename_ack
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_final_index_sum_regn_Sample/$entry
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_final_index_sum_regn_Sample/req
      -- 
    ca_9414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 635_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4455_inst_ack_1, ack => zeropad3D_CP_2152_elements(635)); -- 
    req_9439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(635), ack => array_obj_ref_4461_index_offset_req_0); -- 
    -- CP-element group 636:  transition  input  bypass 
    -- CP-element group 636: predecessors 
    -- CP-element group 636: 	635 
    -- CP-element group 636: successors 
    -- CP-element group 636: 	642 
    -- CP-element group 636:  members (3) 
      -- CP-element group 636: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_final_index_sum_regn_sample_complete
      -- CP-element group 636: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_final_index_sum_regn_Sample/$exit
      -- CP-element group 636: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_final_index_sum_regn_Sample/ack
      -- 
    ack_9440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 636_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4461_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(636)); -- 
    -- CP-element group 637:  transition  input  output  bypass 
    -- CP-element group 637: predecessors 
    -- CP-element group 637: 	1147 
    -- CP-element group 637: successors 
    -- CP-element group 637: 	638 
    -- CP-element group 637:  members (11) 
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/addr_of_4462_sample_start_
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_root_address_calculated
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_offset_calculated
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_final_index_sum_regn_Update/$exit
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_final_index_sum_regn_Update/ack
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_base_plus_offset/$entry
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_base_plus_offset/$exit
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_base_plus_offset/sum_rename_req
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_base_plus_offset/sum_rename_ack
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/addr_of_4462_request/$entry
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/addr_of_4462_request/req
      -- 
    ack_9445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 637_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4461_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(637)); -- 
    req_9454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(637), ack => addr_of_4462_final_reg_req_0); -- 
    -- CP-element group 638:  transition  input  bypass 
    -- CP-element group 638: predecessors 
    -- CP-element group 638: 	637 
    -- CP-element group 638: successors 
    -- CP-element group 638:  members (3) 
      -- CP-element group 638: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/addr_of_4462_sample_completed_
      -- CP-element group 638: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/addr_of_4462_request/$exit
      -- CP-element group 638: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/addr_of_4462_request/ack
      -- 
    ack_9455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 638_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4462_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(638)); -- 
    -- CP-element group 639:  join  fork  transition  input  output  bypass 
    -- CP-element group 639: predecessors 
    -- CP-element group 639: 	1147 
    -- CP-element group 639: successors 
    -- CP-element group 639: 	640 
    -- CP-element group 639:  members (28) 
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/addr_of_4462_update_completed_
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/addr_of_4462_complete/$exit
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/addr_of_4462_complete/ack
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_sample_start_
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_base_address_calculated
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_word_address_calculated
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_root_address_calculated
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_base_address_resized
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_base_addr_resize/$entry
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_base_addr_resize/$exit
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_base_addr_resize/base_resize_req
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_base_addr_resize/base_resize_ack
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_base_plus_offset/$entry
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_base_plus_offset/$exit
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_base_plus_offset/sum_rename_req
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_base_plus_offset/sum_rename_ack
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_word_addrgen/$entry
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_word_addrgen/$exit
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_word_addrgen/root_register_req
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_word_addrgen/root_register_ack
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Sample/$entry
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Sample/ptr_deref_4465_Split/$entry
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Sample/ptr_deref_4465_Split/$exit
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Sample/ptr_deref_4465_Split/split_req
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Sample/ptr_deref_4465_Split/split_ack
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Sample/word_access_start/$entry
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Sample/word_access_start/word_0/$entry
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Sample/word_access_start/word_0/rr
      -- 
    ack_9460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 639_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4462_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(639)); -- 
    rr_9498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(639), ack => ptr_deref_4465_store_0_req_0); -- 
    -- CP-element group 640:  transition  input  bypass 
    -- CP-element group 640: predecessors 
    -- CP-element group 640: 	639 
    -- CP-element group 640: successors 
    -- CP-element group 640:  members (5) 
      -- CP-element group 640: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_sample_completed_
      -- CP-element group 640: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Sample/$exit
      -- CP-element group 640: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Sample/word_access_start/$exit
      -- CP-element group 640: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Sample/word_access_start/word_0/$exit
      -- CP-element group 640: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Sample/word_access_start/word_0/ra
      -- 
    ra_9499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 640_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4465_store_0_ack_0, ack => zeropad3D_CP_2152_elements(640)); -- 
    -- CP-element group 641:  transition  input  bypass 
    -- CP-element group 641: predecessors 
    -- CP-element group 641: 	1147 
    -- CP-element group 641: successors 
    -- CP-element group 641: 	642 
    -- CP-element group 641:  members (5) 
      -- CP-element group 641: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_update_completed_
      -- CP-element group 641: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Update/$exit
      -- CP-element group 641: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Update/word_access_complete/$exit
      -- CP-element group 641: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Update/word_access_complete/word_0/$exit
      -- CP-element group 641: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Update/word_access_complete/word_0/ca
      -- 
    ca_9510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 641_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4465_store_0_ack_1, ack => zeropad3D_CP_2152_elements(641)); -- 
    -- CP-element group 642:  join  transition  place  bypass 
    -- CP-element group 642: predecessors 
    -- CP-element group 642: 	636 
    -- CP-element group 642: 	641 
    -- CP-element group 642: successors 
    -- CP-element group 642: 	1148 
    -- CP-element group 642:  members (5) 
      -- CP-element group 642: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468__exit__
      -- CP-element group 642: 	 branch_block_stmt_714/ifx_xthen1376_ifx_xend1445
      -- CP-element group 642: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/$exit
      -- CP-element group 642: 	 branch_block_stmt_714/ifx_xthen1376_ifx_xend1445_PhiReq/$entry
      -- CP-element group 642: 	 branch_block_stmt_714/ifx_xthen1376_ifx_xend1445_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_642: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_642"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(636) & zeropad3D_CP_2152_elements(641);
      gj_zeropad3D_cp_element_group_642 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(642), clk => clk, reset => reset); --
    end block;
    -- CP-element group 643:  transition  input  bypass 
    -- CP-element group 643: predecessors 
    -- CP-element group 643: 	627 
    -- CP-element group 643: successors 
    -- CP-element group 643:  members (3) 
      -- CP-element group 643: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4474_sample_completed_
      -- CP-element group 643: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4474_Sample/$exit
      -- CP-element group 643: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4474_Sample/ra
      -- 
    ra_9522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 643_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4474_inst_ack_0, ack => zeropad3D_CP_2152_elements(643)); -- 
    -- CP-element group 644:  fork  transition  input  output  bypass 
    -- CP-element group 644: predecessors 
    -- CP-element group 644: 	627 
    -- CP-element group 644: successors 
    -- CP-element group 644: 	645 
    -- CP-element group 644: 	653 
    -- CP-element group 644:  members (9) 
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4474_update_completed_
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4474_Update/$exit
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4474_Update/ca
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4538_sample_start_
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4538_Sample/$entry
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4538_Sample/rr
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4563_sample_start_
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4563_Sample/$entry
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4563_Sample/rr
      -- 
    ca_9527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 644_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4474_inst_ack_1, ack => zeropad3D_CP_2152_elements(644)); -- 
    rr_9535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(644), ack => type_cast_4538_inst_req_0); -- 
    rr_9645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(644), ack => type_cast_4563_inst_req_0); -- 
    -- CP-element group 645:  transition  input  bypass 
    -- CP-element group 645: predecessors 
    -- CP-element group 645: 	644 
    -- CP-element group 645: successors 
    -- CP-element group 645:  members (3) 
      -- CP-element group 645: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4538_sample_completed_
      -- CP-element group 645: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4538_Sample/$exit
      -- CP-element group 645: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4538_Sample/ra
      -- 
    ra_9536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 645_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4538_inst_ack_0, ack => zeropad3D_CP_2152_elements(645)); -- 
    -- CP-element group 646:  transition  input  output  bypass 
    -- CP-element group 646: predecessors 
    -- CP-element group 646: 	627 
    -- CP-element group 646: successors 
    -- CP-element group 646: 	647 
    -- CP-element group 646:  members (16) 
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4538_update_completed_
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4538_Update/$exit
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4538_Update/ca
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_index_resized_1
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_index_scaled_1
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_index_computed_1
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_index_resize_1/$entry
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_index_resize_1/$exit
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_index_resize_1/index_resize_req
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_index_resize_1/index_resize_ack
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_index_scale_1/$entry
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_index_scale_1/$exit
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_index_scale_1/scale_rename_req
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_index_scale_1/scale_rename_ack
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_final_index_sum_regn_Sample/$entry
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_final_index_sum_regn_Sample/req
      -- 
    ca_9541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 646_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4538_inst_ack_1, ack => zeropad3D_CP_2152_elements(646)); -- 
    req_9566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(646), ack => array_obj_ref_4544_index_offset_req_0); -- 
    -- CP-element group 647:  transition  input  bypass 
    -- CP-element group 647: predecessors 
    -- CP-element group 647: 	646 
    -- CP-element group 647: successors 
    -- CP-element group 647: 	662 
    -- CP-element group 647:  members (3) 
      -- CP-element group 647: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_final_index_sum_regn_sample_complete
      -- CP-element group 647: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_final_index_sum_regn_Sample/$exit
      -- CP-element group 647: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_final_index_sum_regn_Sample/ack
      -- 
    ack_9567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 647_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4544_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(647)); -- 
    -- CP-element group 648:  transition  input  output  bypass 
    -- CP-element group 648: predecessors 
    -- CP-element group 648: 	627 
    -- CP-element group 648: successors 
    -- CP-element group 648: 	649 
    -- CP-element group 648:  members (11) 
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4545_sample_start_
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_root_address_calculated
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_offset_calculated
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_final_index_sum_regn_Update/$exit
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_final_index_sum_regn_Update/ack
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_base_plus_offset/$entry
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_base_plus_offset/$exit
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_base_plus_offset/sum_rename_req
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4544_base_plus_offset/sum_rename_ack
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4545_request/$entry
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4545_request/req
      -- 
    ack_9572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 648_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4544_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(648)); -- 
    req_9581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(648), ack => addr_of_4545_final_reg_req_0); -- 
    -- CP-element group 649:  transition  input  bypass 
    -- CP-element group 649: predecessors 
    -- CP-element group 649: 	648 
    -- CP-element group 649: successors 
    -- CP-element group 649:  members (3) 
      -- CP-element group 649: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4545_sample_completed_
      -- CP-element group 649: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4545_request/$exit
      -- CP-element group 649: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4545_request/ack
      -- 
    ack_9582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 649_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4545_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(649)); -- 
    -- CP-element group 650:  join  fork  transition  input  output  bypass 
    -- CP-element group 650: predecessors 
    -- CP-element group 650: 	627 
    -- CP-element group 650: successors 
    -- CP-element group 650: 	651 
    -- CP-element group 650:  members (24) 
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4545_update_completed_
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4545_complete/$exit
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4545_complete/ack
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_sample_start_
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_base_address_calculated
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_word_address_calculated
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_root_address_calculated
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_base_address_resized
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_base_addr_resize/$entry
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_base_addr_resize/$exit
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_base_addr_resize/base_resize_req
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_base_addr_resize/base_resize_ack
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_base_plus_offset/$entry
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_base_plus_offset/$exit
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_base_plus_offset/sum_rename_req
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_base_plus_offset/sum_rename_ack
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_word_addrgen/$entry
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_word_addrgen/$exit
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_word_addrgen/root_register_req
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_word_addrgen/root_register_ack
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Sample/$entry
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Sample/word_access_start/$entry
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Sample/word_access_start/word_0/$entry
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Sample/word_access_start/word_0/rr
      -- 
    ack_9587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 650_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4545_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(650)); -- 
    rr_9620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(650), ack => ptr_deref_4549_load_0_req_0); -- 
    -- CP-element group 651:  transition  input  bypass 
    -- CP-element group 651: predecessors 
    -- CP-element group 651: 	650 
    -- CP-element group 651: successors 
    -- CP-element group 651:  members (5) 
      -- CP-element group 651: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_sample_completed_
      -- CP-element group 651: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Sample/$exit
      -- CP-element group 651: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Sample/word_access_start/$exit
      -- CP-element group 651: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Sample/word_access_start/word_0/$exit
      -- CP-element group 651: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Sample/word_access_start/word_0/ra
      -- 
    ra_9621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 651_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4549_load_0_ack_0, ack => zeropad3D_CP_2152_elements(651)); -- 
    -- CP-element group 652:  transition  input  bypass 
    -- CP-element group 652: predecessors 
    -- CP-element group 652: 	627 
    -- CP-element group 652: successors 
    -- CP-element group 652: 	659 
    -- CP-element group 652:  members (9) 
      -- CP-element group 652: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_update_completed_
      -- CP-element group 652: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Update/$exit
      -- CP-element group 652: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Update/word_access_complete/$exit
      -- CP-element group 652: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Update/word_access_complete/word_0/$exit
      -- CP-element group 652: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Update/word_access_complete/word_0/ca
      -- CP-element group 652: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Update/ptr_deref_4549_Merge/$entry
      -- CP-element group 652: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Update/ptr_deref_4549_Merge/$exit
      -- CP-element group 652: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Update/ptr_deref_4549_Merge/merge_req
      -- CP-element group 652: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4549_Update/ptr_deref_4549_Merge/merge_ack
      -- 
    ca_9632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 652_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4549_load_0_ack_1, ack => zeropad3D_CP_2152_elements(652)); -- 
    -- CP-element group 653:  transition  input  bypass 
    -- CP-element group 653: predecessors 
    -- CP-element group 653: 	644 
    -- CP-element group 653: successors 
    -- CP-element group 653:  members (3) 
      -- CP-element group 653: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4563_sample_completed_
      -- CP-element group 653: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4563_Sample/$exit
      -- CP-element group 653: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4563_Sample/ra
      -- 
    ra_9646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 653_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4563_inst_ack_0, ack => zeropad3D_CP_2152_elements(653)); -- 
    -- CP-element group 654:  transition  input  output  bypass 
    -- CP-element group 654: predecessors 
    -- CP-element group 654: 	627 
    -- CP-element group 654: successors 
    -- CP-element group 654: 	655 
    -- CP-element group 654:  members (16) 
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4563_update_completed_
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4563_Update/$exit
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/type_cast_4563_Update/ca
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_index_resized_1
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_index_scaled_1
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_index_computed_1
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_index_resize_1/$entry
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_index_resize_1/$exit
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_index_resize_1/index_resize_req
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_index_resize_1/index_resize_ack
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_index_scale_1/$entry
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_index_scale_1/$exit
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_index_scale_1/scale_rename_req
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_index_scale_1/scale_rename_ack
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_final_index_sum_regn_Sample/$entry
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_final_index_sum_regn_Sample/req
      -- 
    ca_9651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 654_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4563_inst_ack_1, ack => zeropad3D_CP_2152_elements(654)); -- 
    req_9676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(654), ack => array_obj_ref_4569_index_offset_req_0); -- 
    -- CP-element group 655:  transition  input  bypass 
    -- CP-element group 655: predecessors 
    -- CP-element group 655: 	654 
    -- CP-element group 655: successors 
    -- CP-element group 655: 	662 
    -- CP-element group 655:  members (3) 
      -- CP-element group 655: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_final_index_sum_regn_sample_complete
      -- CP-element group 655: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_final_index_sum_regn_Sample/$exit
      -- CP-element group 655: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_final_index_sum_regn_Sample/ack
      -- 
    ack_9677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 655_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4569_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(655)); -- 
    -- CP-element group 656:  transition  input  output  bypass 
    -- CP-element group 656: predecessors 
    -- CP-element group 656: 	627 
    -- CP-element group 656: successors 
    -- CP-element group 656: 	657 
    -- CP-element group 656:  members (11) 
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4570_sample_start_
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_root_address_calculated
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_offset_calculated
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_final_index_sum_regn_Update/$exit
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_final_index_sum_regn_Update/ack
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_base_plus_offset/$entry
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_base_plus_offset/$exit
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_base_plus_offset/sum_rename_req
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/array_obj_ref_4569_base_plus_offset/sum_rename_ack
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4570_request/$entry
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4570_request/req
      -- 
    ack_9682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 656_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4569_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(656)); -- 
    req_9691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(656), ack => addr_of_4570_final_reg_req_0); -- 
    -- CP-element group 657:  transition  input  bypass 
    -- CP-element group 657: predecessors 
    -- CP-element group 657: 	656 
    -- CP-element group 657: successors 
    -- CP-element group 657:  members (3) 
      -- CP-element group 657: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4570_sample_completed_
      -- CP-element group 657: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4570_request/$exit
      -- CP-element group 657: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4570_request/ack
      -- 
    ack_9692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 657_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4570_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(657)); -- 
    -- CP-element group 658:  fork  transition  input  bypass 
    -- CP-element group 658: predecessors 
    -- CP-element group 658: 	627 
    -- CP-element group 658: successors 
    -- CP-element group 658: 	659 
    -- CP-element group 658:  members (19) 
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4570_update_completed_
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4570_complete/$exit
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/addr_of_4570_complete/ack
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_base_address_calculated
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_word_address_calculated
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_root_address_calculated
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_base_address_resized
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_base_addr_resize/$entry
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_base_addr_resize/$exit
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_base_addr_resize/base_resize_req
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_base_addr_resize/base_resize_ack
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_base_plus_offset/$entry
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_base_plus_offset/$exit
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_base_plus_offset/sum_rename_req
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_base_plus_offset/sum_rename_ack
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_word_addrgen/$entry
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_word_addrgen/$exit
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_word_addrgen/root_register_req
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_word_addrgen/root_register_ack
      -- 
    ack_9697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 658_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4570_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(658)); -- 
    -- CP-element group 659:  join  transition  output  bypass 
    -- CP-element group 659: predecessors 
    -- CP-element group 659: 	652 
    -- CP-element group 659: 	658 
    -- CP-element group 659: successors 
    -- CP-element group 659: 	660 
    -- CP-element group 659:  members (9) 
      -- CP-element group 659: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_sample_start_
      -- CP-element group 659: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Sample/$entry
      -- CP-element group 659: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Sample/ptr_deref_4573_Split/$entry
      -- CP-element group 659: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Sample/ptr_deref_4573_Split/$exit
      -- CP-element group 659: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Sample/ptr_deref_4573_Split/split_req
      -- CP-element group 659: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Sample/ptr_deref_4573_Split/split_ack
      -- CP-element group 659: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Sample/word_access_start/$entry
      -- CP-element group 659: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Sample/word_access_start/word_0/$entry
      -- CP-element group 659: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Sample/word_access_start/word_0/rr
      -- 
    rr_9735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(659), ack => ptr_deref_4573_store_0_req_0); -- 
    zeropad3D_cp_element_group_659: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_659"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(652) & zeropad3D_CP_2152_elements(658);
      gj_zeropad3D_cp_element_group_659 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(659), clk => clk, reset => reset); --
    end block;
    -- CP-element group 660:  transition  input  bypass 
    -- CP-element group 660: predecessors 
    -- CP-element group 660: 	659 
    -- CP-element group 660: successors 
    -- CP-element group 660:  members (5) 
      -- CP-element group 660: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_sample_completed_
      -- CP-element group 660: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Sample/$exit
      -- CP-element group 660: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Sample/word_access_start/$exit
      -- CP-element group 660: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Sample/word_access_start/word_0/$exit
      -- CP-element group 660: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Sample/word_access_start/word_0/ra
      -- 
    ra_9736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 660_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4573_store_0_ack_0, ack => zeropad3D_CP_2152_elements(660)); -- 
    -- CP-element group 661:  transition  input  bypass 
    -- CP-element group 661: predecessors 
    -- CP-element group 661: 	627 
    -- CP-element group 661: successors 
    -- CP-element group 661: 	662 
    -- CP-element group 661:  members (5) 
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Update/word_access_complete/word_0/ca
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Update/word_access_complete/$exit
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Update/word_access_complete/word_0/$exit
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_update_completed_
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/ptr_deref_4573_Update/$exit
      -- 
    ca_9747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 661_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4573_store_0_ack_1, ack => zeropad3D_CP_2152_elements(661)); -- 
    -- CP-element group 662:  join  transition  place  bypass 
    -- CP-element group 662: predecessors 
    -- CP-element group 662: 	647 
    -- CP-element group 662: 	655 
    -- CP-element group 662: 	661 
    -- CP-element group 662: successors 
    -- CP-element group 662: 	1148 
    -- CP-element group 662:  members (5) 
      -- CP-element group 662: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575__exit__
      -- CP-element group 662: 	 branch_block_stmt_714/ifx_xelse1397_ifx_xend1445
      -- CP-element group 662: 	 branch_block_stmt_714/assign_stmt_4475_to_assign_stmt_4575/$exit
      -- CP-element group 662: 	 branch_block_stmt_714/ifx_xelse1397_ifx_xend1445_PhiReq/$entry
      -- CP-element group 662: 	 branch_block_stmt_714/ifx_xelse1397_ifx_xend1445_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_662: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_662"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(647) & zeropad3D_CP_2152_elements(655) & zeropad3D_CP_2152_elements(661);
      gj_zeropad3D_cp_element_group_662 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(662), clk => clk, reset => reset); --
    end block;
    -- CP-element group 663:  transition  input  bypass 
    -- CP-element group 663: predecessors 
    -- CP-element group 663: 	1148 
    -- CP-element group 663: successors 
    -- CP-element group 663:  members (3) 
      -- CP-element group 663: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/type_cast_4581_sample_completed_
      -- CP-element group 663: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/type_cast_4581_Sample/ra
      -- CP-element group 663: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/type_cast_4581_Sample/$exit
      -- 
    ra_9759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 663_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4581_inst_ack_0, ack => zeropad3D_CP_2152_elements(663)); -- 
    -- CP-element group 664:  branch  transition  place  input  output  bypass 
    -- CP-element group 664: predecessors 
    -- CP-element group 664: 	1148 
    -- CP-element group 664: successors 
    -- CP-element group 664: 	665 
    -- CP-element group 664: 	666 
    -- CP-element group 664:  members (13) 
      -- CP-element group 664: 	 branch_block_stmt_714/if_stmt_4596__entry__
      -- CP-element group 664: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595__exit__
      -- CP-element group 664: 	 branch_block_stmt_714/if_stmt_4596_else_link/$entry
      -- CP-element group 664: 	 branch_block_stmt_714/if_stmt_4596_if_link/$entry
      -- CP-element group 664: 	 branch_block_stmt_714/if_stmt_4596_eval_test/branch_req
      -- CP-element group 664: 	 branch_block_stmt_714/if_stmt_4596_eval_test/$exit
      -- CP-element group 664: 	 branch_block_stmt_714/if_stmt_4596_eval_test/$entry
      -- CP-element group 664: 	 branch_block_stmt_714/if_stmt_4596_dead_link/$entry
      -- CP-element group 664: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/type_cast_4581_Update/ca
      -- CP-element group 664: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/$exit
      -- CP-element group 664: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/type_cast_4581_Update/$exit
      -- CP-element group 664: 	 branch_block_stmt_714/R_cmp1453_4597_place
      -- CP-element group 664: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/type_cast_4581_update_completed_
      -- 
    ca_9764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 664_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4581_inst_ack_1, ack => zeropad3D_CP_2152_elements(664)); -- 
    branch_req_9772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(664), ack => if_stmt_4596_branch_req_0); -- 
    -- CP-element group 665:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 665: predecessors 
    -- CP-element group 665: 	664 
    -- CP-element group 665: successors 
    -- CP-element group 665: 	1157 
    -- CP-element group 665: 	1158 
    -- CP-element group 665: 	1160 
    -- CP-element group 665: 	1161 
    -- CP-element group 665: 	1163 
    -- CP-element group 665: 	1164 
    -- CP-element group 665:  members (40) 
      -- CP-element group 665: 	 branch_block_stmt_714/assign_stmt_4608__entry__
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496
      -- CP-element group 665: 	 branch_block_stmt_714/merge_stmt_4602__exit__
      -- CP-element group 665: 	 branch_block_stmt_714/assign_stmt_4608__exit__
      -- CP-element group 665: 	 branch_block_stmt_714/assign_stmt_4608/$exit
      -- CP-element group 665: 	 branch_block_stmt_714/assign_stmt_4608/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/if_stmt_4596_if_link/if_choice_transition
      -- CP-element group 665: 	 branch_block_stmt_714/if_stmt_4596_if_link/$exit
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xend1445_ifx_xthen1455
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xend1445_ifx_xthen1455_PhiReq/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xend1445_ifx_xthen1455_PhiReq/$exit
      -- CP-element group 665: 	 branch_block_stmt_714/merge_stmt_4602_PhiReqMerge
      -- CP-element group 665: 	 branch_block_stmt_714/merge_stmt_4602_PhiAck/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/merge_stmt_4602_PhiAck/$exit
      -- CP-element group 665: 	 branch_block_stmt_714/merge_stmt_4602_PhiAck/dummy
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4708/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4708/SplitProtocol/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4708/SplitProtocol/Sample/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4708/SplitProtocol/Sample/rr
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4708/SplitProtocol/Update/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4708/SplitProtocol/Update/cr
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4700/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4700/SplitProtocol/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4700/SplitProtocol/Sample/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4700/SplitProtocol/Sample/rr
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4700/SplitProtocol/Update/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4700/SplitProtocol/Update/cr
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/type_cast_4696/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/type_cast_4696/SplitProtocol/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/type_cast_4696/SplitProtocol/Sample/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/type_cast_4696/SplitProtocol/Sample/rr
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/type_cast_4696/SplitProtocol/Update/$entry
      -- CP-element group 665: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/type_cast_4696/SplitProtocol/Update/cr
      -- 
    if_choice_transition_9777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 665_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4596_branch_ack_1, ack => zeropad3D_CP_2152_elements(665)); -- 
    rr_13803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(665), ack => type_cast_4708_inst_req_0); -- 
    cr_13808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(665), ack => type_cast_4708_inst_req_1); -- 
    rr_13826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(665), ack => type_cast_4700_inst_req_0); -- 
    cr_13831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(665), ack => type_cast_4700_inst_req_1); -- 
    rr_13849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(665), ack => type_cast_4696_inst_req_0); -- 
    cr_13854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(665), ack => type_cast_4696_inst_req_1); -- 
    -- CP-element group 666:  fork  transition  place  input  output  bypass 
    -- CP-element group 666: predecessors 
    -- CP-element group 666: 	664 
    -- CP-element group 666: successors 
    -- CP-element group 666: 	667 
    -- CP-element group 666: 	668 
    -- CP-element group 666: 	669 
    -- CP-element group 666: 	670 
    -- CP-element group 666: 	672 
    -- CP-element group 666: 	675 
    -- CP-element group 666: 	677 
    -- CP-element group 666: 	678 
    -- CP-element group 666: 	679 
    -- CP-element group 666: 	681 
    -- CP-element group 666:  members (54) 
      -- CP-element group 666: 	 branch_block_stmt_714/merge_stmt_4610__exit__
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682__entry__
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4620_Sample/rr
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_update_start_
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4664_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4664_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_word_address_calculated
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_sample_start_
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4620_Sample/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4620_update_start_
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4620_sample_start_
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/if_stmt_4596_else_link/else_choice_transition
      -- CP-element group 666: 	 branch_block_stmt_714/if_stmt_4596_else_link/$exit
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Sample/word_access_start/word_0/rr
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4664_update_start_
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Update/word_access_complete/word_0/cr
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4647_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Update/word_access_complete/word_0/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Sample/word_access_start/word_0/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Update/word_access_complete/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/ifx_xend1445_ifx_xelse1460
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4647_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_sample_start_
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Sample/word_access_start/word_0/rr
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4647_update_start_
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Sample/word_access_start/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Sample/word_access_start/word_0/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4627_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4627_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Sample/word_access_start/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4627_update_start_
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4620_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Sample/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_root_address_calculated
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Sample/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_word_address_calculated
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_root_address_calculated
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Update/word_access_complete/word_0/cr
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4671_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4620_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_update_start_
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Update/word_access_complete/word_0/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Update/word_access_complete/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4671_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4671_update_start_
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/ifx_xend1445_ifx_xelse1460_PhiReq/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/ifx_xend1445_ifx_xelse1460_PhiReq/$exit
      -- CP-element group 666: 	 branch_block_stmt_714/merge_stmt_4610_PhiReqMerge
      -- CP-element group 666: 	 branch_block_stmt_714/merge_stmt_4610_PhiAck/$entry
      -- CP-element group 666: 	 branch_block_stmt_714/merge_stmt_4610_PhiAck/$exit
      -- CP-element group 666: 	 branch_block_stmt_714/merge_stmt_4610_PhiAck/dummy
      -- 
    else_choice_transition_9781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 666_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4596_branch_ack_0, ack => zeropad3D_CP_2152_elements(666)); -- 
    rr_9797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(666), ack => type_cast_4620_inst_req_0); -- 
    cr_9877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(666), ack => type_cast_4664_inst_req_1); -- 
    rr_9819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(666), ack => LOAD_col_high_4623_load_0_req_0); -- 
    cr_9905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(666), ack => LOAD_row_high_4667_load_0_req_1); -- 
    cr_9863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(666), ack => type_cast_4647_inst_req_1); -- 
    rr_9894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(666), ack => LOAD_row_high_4667_load_0_req_0); -- 
    cr_9849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(666), ack => type_cast_4627_inst_req_1); -- 
    cr_9802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(666), ack => type_cast_4620_inst_req_1); -- 
    cr_9830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(666), ack => LOAD_col_high_4623_load_0_req_1); -- 
    cr_9924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(666), ack => type_cast_4671_inst_req_1); -- 
    -- CP-element group 667:  transition  input  bypass 
    -- CP-element group 667: predecessors 
    -- CP-element group 667: 	666 
    -- CP-element group 667: successors 
    -- CP-element group 667:  members (3) 
      -- CP-element group 667: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4620_Sample/$exit
      -- CP-element group 667: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4620_sample_completed_
      -- CP-element group 667: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4620_Sample/ra
      -- 
    ra_9798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 667_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4620_inst_ack_0, ack => zeropad3D_CP_2152_elements(667)); -- 
    -- CP-element group 668:  transition  input  bypass 
    -- CP-element group 668: predecessors 
    -- CP-element group 668: 	666 
    -- CP-element group 668: successors 
    -- CP-element group 668: 	673 
    -- CP-element group 668:  members (3) 
      -- CP-element group 668: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4620_update_completed_
      -- CP-element group 668: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4620_Update/ca
      -- CP-element group 668: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4620_Update/$exit
      -- 
    ca_9803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 668_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4620_inst_ack_1, ack => zeropad3D_CP_2152_elements(668)); -- 
    -- CP-element group 669:  transition  input  bypass 
    -- CP-element group 669: predecessors 
    -- CP-element group 669: 	666 
    -- CP-element group 669: successors 
    -- CP-element group 669:  members (5) 
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Sample/word_access_start/word_0/ra
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Sample/word_access_start/word_0/$exit
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_sample_completed_
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Sample/word_access_start/$exit
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Sample/$exit
      -- 
    ra_9820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 669_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4623_load_0_ack_0, ack => zeropad3D_CP_2152_elements(669)); -- 
    -- CP-element group 670:  transition  input  output  bypass 
    -- CP-element group 670: predecessors 
    -- CP-element group 670: 	666 
    -- CP-element group 670: successors 
    -- CP-element group 670: 	671 
    -- CP-element group 670:  members (12) 
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_update_completed_
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4627_Sample/rr
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4627_Sample/$entry
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4627_sample_start_
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Update/LOAD_col_high_4623_Merge/merge_ack
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Update/LOAD_col_high_4623_Merge/merge_req
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Update/LOAD_col_high_4623_Merge/$exit
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Update/LOAD_col_high_4623_Merge/$entry
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Update/word_access_complete/word_0/ca
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Update/word_access_complete/word_0/$exit
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Update/word_access_complete/$exit
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_col_high_4623_Update/$exit
      -- 
    ca_9831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 670_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4623_load_0_ack_1, ack => zeropad3D_CP_2152_elements(670)); -- 
    rr_9844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(670), ack => type_cast_4627_inst_req_0); -- 
    -- CP-element group 671:  transition  input  bypass 
    -- CP-element group 671: predecessors 
    -- CP-element group 671: 	670 
    -- CP-element group 671: successors 
    -- CP-element group 671:  members (3) 
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4627_Sample/ra
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4627_Sample/$exit
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4627_sample_completed_
      -- 
    ra_9845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 671_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4627_inst_ack_0, ack => zeropad3D_CP_2152_elements(671)); -- 
    -- CP-element group 672:  transition  input  bypass 
    -- CP-element group 672: predecessors 
    -- CP-element group 672: 	666 
    -- CP-element group 672: successors 
    -- CP-element group 672: 	673 
    -- CP-element group 672:  members (3) 
      -- CP-element group 672: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4627_Update/ca
      -- CP-element group 672: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4627_Update/$exit
      -- CP-element group 672: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4627_update_completed_
      -- 
    ca_9850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 672_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4627_inst_ack_1, ack => zeropad3D_CP_2152_elements(672)); -- 
    -- CP-element group 673:  join  transition  output  bypass 
    -- CP-element group 673: predecessors 
    -- CP-element group 673: 	668 
    -- CP-element group 673: 	672 
    -- CP-element group 673: successors 
    -- CP-element group 673: 	674 
    -- CP-element group 673:  members (3) 
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4647_Sample/rr
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4647_Sample/$entry
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4647_sample_start_
      -- 
    rr_9858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(673), ack => type_cast_4647_inst_req_0); -- 
    zeropad3D_cp_element_group_673: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_673"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(668) & zeropad3D_CP_2152_elements(672);
      gj_zeropad3D_cp_element_group_673 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(673), clk => clk, reset => reset); --
    end block;
    -- CP-element group 674:  transition  input  bypass 
    -- CP-element group 674: predecessors 
    -- CP-element group 674: 	673 
    -- CP-element group 674: successors 
    -- CP-element group 674:  members (3) 
      -- CP-element group 674: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4647_Sample/ra
      -- CP-element group 674: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4647_Sample/$exit
      -- CP-element group 674: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4647_sample_completed_
      -- 
    ra_9859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 674_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4647_inst_ack_0, ack => zeropad3D_CP_2152_elements(674)); -- 
    -- CP-element group 675:  transition  input  output  bypass 
    -- CP-element group 675: predecessors 
    -- CP-element group 675: 	666 
    -- CP-element group 675: successors 
    -- CP-element group 675: 	676 
    -- CP-element group 675:  members (6) 
      -- CP-element group 675: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4664_Sample/rr
      -- CP-element group 675: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4664_Sample/$entry
      -- CP-element group 675: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4664_sample_start_
      -- CP-element group 675: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4647_Update/ca
      -- CP-element group 675: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4647_Update/$exit
      -- CP-element group 675: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4647_update_completed_
      -- 
    ca_9864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 675_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4647_inst_ack_1, ack => zeropad3D_CP_2152_elements(675)); -- 
    rr_9872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(675), ack => type_cast_4664_inst_req_0); -- 
    -- CP-element group 676:  transition  input  bypass 
    -- CP-element group 676: predecessors 
    -- CP-element group 676: 	675 
    -- CP-element group 676: successors 
    -- CP-element group 676:  members (3) 
      -- CP-element group 676: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4664_Sample/ra
      -- CP-element group 676: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4664_Sample/$exit
      -- CP-element group 676: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4664_sample_completed_
      -- 
    ra_9873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 676_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4664_inst_ack_0, ack => zeropad3D_CP_2152_elements(676)); -- 
    -- CP-element group 677:  transition  input  bypass 
    -- CP-element group 677: predecessors 
    -- CP-element group 677: 	666 
    -- CP-element group 677: successors 
    -- CP-element group 677: 	682 
    -- CP-element group 677:  members (3) 
      -- CP-element group 677: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4664_Update/$exit
      -- CP-element group 677: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4664_Update/ca
      -- CP-element group 677: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4664_update_completed_
      -- 
    ca_9878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 677_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4664_inst_ack_1, ack => zeropad3D_CP_2152_elements(677)); -- 
    -- CP-element group 678:  transition  input  bypass 
    -- CP-element group 678: predecessors 
    -- CP-element group 678: 	666 
    -- CP-element group 678: successors 
    -- CP-element group 678:  members (5) 
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Sample/word_access_start/word_0/ra
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Sample/word_access_start/word_0/$exit
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Sample/word_access_start/$exit
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Sample/$exit
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_sample_completed_
      -- 
    ra_9895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 678_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4667_load_0_ack_0, ack => zeropad3D_CP_2152_elements(678)); -- 
    -- CP-element group 679:  transition  input  output  bypass 
    -- CP-element group 679: predecessors 
    -- CP-element group 679: 	666 
    -- CP-element group 679: successors 
    -- CP-element group 679: 	680 
    -- CP-element group 679:  members (12) 
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4671_sample_start_
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Update/LOAD_row_high_4667_Merge/merge_ack
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Update/LOAD_row_high_4667_Merge/merge_req
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Update/LOAD_row_high_4667_Merge/$exit
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Update/LOAD_row_high_4667_Merge/$entry
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Update/word_access_complete/word_0/ca
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Update/word_access_complete/word_0/$exit
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Update/word_access_complete/$exit
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_Update/$exit
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/LOAD_row_high_4667_update_completed_
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4671_Sample/rr
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4671_Sample/$entry
      -- 
    ca_9906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 679_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4667_load_0_ack_1, ack => zeropad3D_CP_2152_elements(679)); -- 
    rr_9919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(679), ack => type_cast_4671_inst_req_0); -- 
    -- CP-element group 680:  transition  input  bypass 
    -- CP-element group 680: predecessors 
    -- CP-element group 680: 	679 
    -- CP-element group 680: successors 
    -- CP-element group 680:  members (3) 
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4671_Sample/ra
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4671_Sample/$exit
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4671_sample_completed_
      -- 
    ra_9920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 680_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4671_inst_ack_0, ack => zeropad3D_CP_2152_elements(680)); -- 
    -- CP-element group 681:  transition  input  bypass 
    -- CP-element group 681: predecessors 
    -- CP-element group 681: 	666 
    -- CP-element group 681: successors 
    -- CP-element group 681: 	682 
    -- CP-element group 681:  members (3) 
      -- CP-element group 681: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4671_Update/ca
      -- CP-element group 681: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4671_Update/$exit
      -- CP-element group 681: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/type_cast_4671_update_completed_
      -- 
    ca_9925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 681_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4671_inst_ack_1, ack => zeropad3D_CP_2152_elements(681)); -- 
    -- CP-element group 682:  branch  join  transition  place  output  bypass 
    -- CP-element group 682: predecessors 
    -- CP-element group 682: 	677 
    -- CP-element group 682: 	681 
    -- CP-element group 682: successors 
    -- CP-element group 682: 	683 
    -- CP-element group 682: 	684 
    -- CP-element group 682:  members (10) 
      -- CP-element group 682: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682__exit__
      -- CP-element group 682: 	 branch_block_stmt_714/if_stmt_4683__entry__
      -- CP-element group 682: 	 branch_block_stmt_714/assign_stmt_4616_to_assign_stmt_4682/$exit
      -- CP-element group 682: 	 branch_block_stmt_714/R_cmp1487_4684_place
      -- CP-element group 682: 	 branch_block_stmt_714/if_stmt_4683_else_link/$entry
      -- CP-element group 682: 	 branch_block_stmt_714/if_stmt_4683_if_link/$entry
      -- CP-element group 682: 	 branch_block_stmt_714/if_stmt_4683_eval_test/branch_req
      -- CP-element group 682: 	 branch_block_stmt_714/if_stmt_4683_eval_test/$exit
      -- CP-element group 682: 	 branch_block_stmt_714/if_stmt_4683_eval_test/$entry
      -- CP-element group 682: 	 branch_block_stmt_714/if_stmt_4683_dead_link/$entry
      -- 
    branch_req_9933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(682), ack => if_stmt_4683_branch_req_0); -- 
    zeropad3D_cp_element_group_682: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_682"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(677) & zeropad3D_CP_2152_elements(681);
      gj_zeropad3D_cp_element_group_682 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(682), clk => clk, reset => reset); --
    end block;
    -- CP-element group 683:  fork  transition  place  input  output  bypass 
    -- CP-element group 683: predecessors 
    -- CP-element group 683: 	682 
    -- CP-element group 683: successors 
    -- CP-element group 683: 	1172 
    -- CP-element group 683: 	1173 
    -- CP-element group 683: 	1175 
    -- CP-element group 683: 	1176 
    -- CP-element group 683: 	1178 
    -- CP-element group 683: 	1179 
    -- CP-element group 683:  members (28) 
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497
      -- CP-element group 683: 	 branch_block_stmt_714/if_stmt_4683_if_link/if_choice_transition
      -- CP-element group 683: 	 branch_block_stmt_714/if_stmt_4683_if_link/$exit
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/type_cast_4719/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/type_cast_4719/SplitProtocol/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/type_cast_4719/SplitProtocol/Sample/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/type_cast_4719/SplitProtocol/Sample/rr
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/type_cast_4719/SplitProtocol/Update/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/type_cast_4719/SplitProtocol/Update/cr
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/type_cast_4715/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/type_cast_4715/SplitProtocol/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/type_cast_4715/SplitProtocol/Sample/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/type_cast_4715/SplitProtocol/Sample/rr
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/type_cast_4715/SplitProtocol/Update/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/type_cast_4715/SplitProtocol/Update/cr
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/type_cast_4723/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/type_cast_4723/SplitProtocol/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/type_cast_4723/SplitProtocol/Sample/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/type_cast_4723/SplitProtocol/Sample/rr
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/type_cast_4723/SplitProtocol/Update/$entry
      -- CP-element group 683: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/type_cast_4723/SplitProtocol/Update/cr
      -- 
    if_choice_transition_9938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 683_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4683_branch_ack_1, ack => zeropad3D_CP_2152_elements(683)); -- 
    rr_13882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(683), ack => type_cast_4719_inst_req_0); -- 
    cr_13887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(683), ack => type_cast_4719_inst_req_1); -- 
    rr_13905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(683), ack => type_cast_4715_inst_req_0); -- 
    cr_13910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(683), ack => type_cast_4715_inst_req_1); -- 
    rr_13928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(683), ack => type_cast_4723_inst_req_0); -- 
    cr_13933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(683), ack => type_cast_4723_inst_req_1); -- 
    -- CP-element group 684:  fork  transition  place  input  output  bypass 
    -- CP-element group 684: predecessors 
    -- CP-element group 684: 	682 
    -- CP-element group 684: successors 
    -- CP-element group 684: 	1149 
    -- CP-element group 684: 	1150 
    -- CP-element group 684: 	1152 
    -- CP-element group 684: 	1153 
    -- CP-element group 684: 	1155 
    -- CP-element group 684:  members (22) 
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496
      -- CP-element group 684: 	 branch_block_stmt_714/if_stmt_4683_else_link/else_choice_transition
      -- CP-element group 684: 	 branch_block_stmt_714/if_stmt_4683_else_link/$exit
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4706/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4706/SplitProtocol/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4706/SplitProtocol/Sample/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4706/SplitProtocol/Sample/rr
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4706/SplitProtocol/Update/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4706/SplitProtocol/Update/cr
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4702/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4702/SplitProtocol/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4702/SplitProtocol/Sample/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4702/SplitProtocol/Sample/rr
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4702/SplitProtocol/Update/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4702/SplitProtocol/Update/cr
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4690/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/$entry
      -- 
    else_choice_transition_9942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 684_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4683_branch_ack_0, ack => zeropad3D_CP_2152_elements(684)); -- 
    rr_13746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(684), ack => type_cast_4706_inst_req_0); -- 
    cr_13751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(684), ack => type_cast_4706_inst_req_1); -- 
    rr_13769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(684), ack => type_cast_4702_inst_req_0); -- 
    cr_13774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(684), ack => type_cast_4702_inst_req_1); -- 
    -- CP-element group 685:  transition  input  bypass 
    -- CP-element group 685: predecessors 
    -- CP-element group 685: 	1185 
    -- CP-element group 685: successors 
    -- CP-element group 685:  members (3) 
      -- CP-element group 685: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4727_Sample/ra
      -- CP-element group 685: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4727_Sample/$exit
      -- CP-element group 685: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4727_sample_completed_
      -- 
    ra_9956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 685_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4727_inst_ack_0, ack => zeropad3D_CP_2152_elements(685)); -- 
    -- CP-element group 686:  transition  input  bypass 
    -- CP-element group 686: predecessors 
    -- CP-element group 686: 	1185 
    -- CP-element group 686: successors 
    -- CP-element group 686: 	701 
    -- CP-element group 686:  members (3) 
      -- CP-element group 686: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4727_Update/ca
      -- CP-element group 686: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4727_Update/$exit
      -- CP-element group 686: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4727_update_completed_
      -- 
    ca_9961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 686_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4727_inst_ack_1, ack => zeropad3D_CP_2152_elements(686)); -- 
    -- CP-element group 687:  transition  input  bypass 
    -- CP-element group 687: predecessors 
    -- CP-element group 687: 	1185 
    -- CP-element group 687: successors 
    -- CP-element group 687:  members (3) 
      -- CP-element group 687: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4737_Sample/ra
      -- CP-element group 687: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4737_Sample/$exit
      -- CP-element group 687: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4737_sample_completed_
      -- 
    ra_9970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 687_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4737_inst_ack_0, ack => zeropad3D_CP_2152_elements(687)); -- 
    -- CP-element group 688:  transition  input  bypass 
    -- CP-element group 688: predecessors 
    -- CP-element group 688: 	1185 
    -- CP-element group 688: successors 
    -- CP-element group 688: 	701 
    -- CP-element group 688:  members (3) 
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4737_Update/ca
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4737_Update/$exit
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4737_update_completed_
      -- 
    ca_9975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 688_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4737_inst_ack_1, ack => zeropad3D_CP_2152_elements(688)); -- 
    -- CP-element group 689:  transition  input  bypass 
    -- CP-element group 689: predecessors 
    -- CP-element group 689: 	1185 
    -- CP-element group 689: successors 
    -- CP-element group 689:  members (5) 
      -- CP-element group 689: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Sample/$exit
      -- CP-element group 689: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Sample/word_access_start/$exit
      -- CP-element group 689: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_sample_completed_
      -- CP-element group 689: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Sample/word_access_start/word_0/ra
      -- CP-element group 689: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Sample/word_access_start/word_0/$exit
      -- 
    ra_9992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 689_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_4752_load_0_ack_0, ack => zeropad3D_CP_2152_elements(689)); -- 
    -- CP-element group 690:  transition  input  output  bypass 
    -- CP-element group 690: predecessors 
    -- CP-element group 690: 	1185 
    -- CP-element group 690: successors 
    -- CP-element group 690: 	699 
    -- CP-element group 690:  members (12) 
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4822_sample_start_
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4822_Sample/rr
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_update_completed_
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4822_Sample/$entry
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Update/LOAD_pad_4752_Merge/merge_ack
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Update/LOAD_pad_4752_Merge/merge_req
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Update/LOAD_pad_4752_Merge/$exit
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Update/LOAD_pad_4752_Merge/$entry
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Update/word_access_complete/word_0/ca
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Update/word_access_complete/word_0/$exit
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Update/word_access_complete/$exit
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Update/$exit
      -- 
    ca_10003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 690_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_4752_load_0_ack_1, ack => zeropad3D_CP_2152_elements(690)); -- 
    rr_10163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(690), ack => type_cast_4822_inst_req_0); -- 
    -- CP-element group 691:  transition  input  bypass 
    -- CP-element group 691: predecessors 
    -- CP-element group 691: 	1185 
    -- CP-element group 691: successors 
    -- CP-element group 691:  members (5) 
      -- CP-element group 691: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Sample/word_access_start/word_0/ra
      -- CP-element group 691: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Sample/word_access_start/word_0/$exit
      -- CP-element group 691: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Sample/word_access_start/$exit
      -- CP-element group 691: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Sample/$exit
      -- CP-element group 691: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_sample_completed_
      -- 
    ra_10025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 691_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_4755_load_0_ack_0, ack => zeropad3D_CP_2152_elements(691)); -- 
    -- CP-element group 692:  transition  input  output  bypass 
    -- CP-element group 692: predecessors 
    -- CP-element group 692: 	1185 
    -- CP-element group 692: successors 
    -- CP-element group 692: 	697 
    -- CP-element group 692:  members (12) 
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4783_Sample/rr
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Update/LOAD_depth_high_4755_Merge/merge_ack
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4783_Sample/$entry
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Update/LOAD_depth_high_4755_Merge/merge_req
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Update/LOAD_depth_high_4755_Merge/$exit
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Update/LOAD_depth_high_4755_Merge/$entry
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Update/word_access_complete/word_0/ca
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Update/word_access_complete/word_0/$exit
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Update/word_access_complete/$exit
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4783_sample_start_
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Update/$exit
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_update_completed_
      -- 
    ca_10036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 692_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_4755_load_0_ack_1, ack => zeropad3D_CP_2152_elements(692)); -- 
    rr_10149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(692), ack => type_cast_4783_inst_req_0); -- 
    -- CP-element group 693:  transition  input  bypass 
    -- CP-element group 693: predecessors 
    -- CP-element group 693: 	1185 
    -- CP-element group 693: successors 
    -- CP-element group 693:  members (5) 
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_sample_completed_
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Sample/word_access_start/word_0/ra
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Sample/word_access_start/word_0/$exit
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Sample/word_access_start/$exit
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Sample/$exit
      -- 
    ra_10075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 693_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4767_load_0_ack_0, ack => zeropad3D_CP_2152_elements(693)); -- 
    -- CP-element group 694:  transition  input  bypass 
    -- CP-element group 694: predecessors 
    -- CP-element group 694: 	1185 
    -- CP-element group 694: successors 
    -- CP-element group 694: 	701 
    -- CP-element group 694:  members (9) 
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_update_completed_
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Update/ptr_deref_4767_Merge/merge_ack
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Update/ptr_deref_4767_Merge/merge_req
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Update/ptr_deref_4767_Merge/$exit
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Update/ptr_deref_4767_Merge/$entry
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Update/word_access_complete/word_0/ca
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Update/word_access_complete/word_0/$exit
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Update/word_access_complete/$exit
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Update/$exit
      -- 
    ca_10086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 694_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4767_load_0_ack_1, ack => zeropad3D_CP_2152_elements(694)); -- 
    -- CP-element group 695:  transition  input  bypass 
    -- CP-element group 695: predecessors 
    -- CP-element group 695: 	1185 
    -- CP-element group 695: successors 
    -- CP-element group 695:  members (5) 
      -- CP-element group 695: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Sample/word_access_start/word_0/ra
      -- CP-element group 695: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_sample_completed_
      -- CP-element group 695: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Sample/word_access_start/word_0/$exit
      -- CP-element group 695: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Sample/word_access_start/$exit
      -- CP-element group 695: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Sample/$exit
      -- 
    ra_10125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 695_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4779_load_0_ack_0, ack => zeropad3D_CP_2152_elements(695)); -- 
    -- CP-element group 696:  transition  input  bypass 
    -- CP-element group 696: predecessors 
    -- CP-element group 696: 	1185 
    -- CP-element group 696: successors 
    -- CP-element group 696: 	701 
    -- CP-element group 696:  members (9) 
      -- CP-element group 696: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Update/$exit
      -- CP-element group 696: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_update_completed_
      -- CP-element group 696: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Update/ptr_deref_4779_Merge/merge_ack
      -- CP-element group 696: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Update/ptr_deref_4779_Merge/merge_req
      -- CP-element group 696: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Update/ptr_deref_4779_Merge/$exit
      -- CP-element group 696: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Update/ptr_deref_4779_Merge/$entry
      -- CP-element group 696: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Update/word_access_complete/word_0/ca
      -- CP-element group 696: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Update/word_access_complete/word_0/$exit
      -- CP-element group 696: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Update/word_access_complete/$exit
      -- 
    ca_10136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 696_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4779_load_0_ack_1, ack => zeropad3D_CP_2152_elements(696)); -- 
    -- CP-element group 697:  transition  input  bypass 
    -- CP-element group 697: predecessors 
    -- CP-element group 697: 	692 
    -- CP-element group 697: successors 
    -- CP-element group 697:  members (3) 
      -- CP-element group 697: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4783_Sample/ra
      -- CP-element group 697: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4783_Sample/$exit
      -- CP-element group 697: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4783_sample_completed_
      -- 
    ra_10150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 697_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4783_inst_ack_0, ack => zeropad3D_CP_2152_elements(697)); -- 
    -- CP-element group 698:  transition  input  bypass 
    -- CP-element group 698: predecessors 
    -- CP-element group 698: 	1185 
    -- CP-element group 698: successors 
    -- CP-element group 698: 	701 
    -- CP-element group 698:  members (3) 
      -- CP-element group 698: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4783_Update/ca
      -- CP-element group 698: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4783_Update/$exit
      -- CP-element group 698: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4783_update_completed_
      -- 
    ca_10155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 698_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4783_inst_ack_1, ack => zeropad3D_CP_2152_elements(698)); -- 
    -- CP-element group 699:  transition  input  bypass 
    -- CP-element group 699: predecessors 
    -- CP-element group 699: 	690 
    -- CP-element group 699: successors 
    -- CP-element group 699:  members (3) 
      -- CP-element group 699: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4822_Sample/ra
      -- CP-element group 699: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4822_Sample/$exit
      -- CP-element group 699: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4822_sample_completed_
      -- 
    ra_10164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 699_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4822_inst_ack_0, ack => zeropad3D_CP_2152_elements(699)); -- 
    -- CP-element group 700:  transition  input  bypass 
    -- CP-element group 700: predecessors 
    -- CP-element group 700: 	1185 
    -- CP-element group 700: successors 
    -- CP-element group 700: 	701 
    -- CP-element group 700:  members (3) 
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4822_update_completed_
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4822_Update/$exit
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4822_Update/ca
      -- 
    ca_10169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 700_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4822_inst_ack_1, ack => zeropad3D_CP_2152_elements(700)); -- 
    -- CP-element group 701:  join  fork  transition  place  output  bypass 
    -- CP-element group 701: predecessors 
    -- CP-element group 701: 	686 
    -- CP-element group 701: 	688 
    -- CP-element group 701: 	694 
    -- CP-element group 701: 	696 
    -- CP-element group 701: 	698 
    -- CP-element group 701: 	700 
    -- CP-element group 701: successors 
    -- CP-element group 701: 	1196 
    -- CP-element group 701: 	1197 
    -- CP-element group 701: 	1199 
    -- CP-element group 701: 	1200 
    -- CP-element group 701: 	1202 
    -- CP-element group 701:  members (22) 
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562
      -- CP-element group 701: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864__exit__
      -- CP-element group 701: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/$exit
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4877/SplitProtocol/Sample/rr
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4867/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4885/SplitProtocol/Update/cr
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4885/SplitProtocol/Update/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4885/SplitProtocol/Sample/rr
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4885/SplitProtocol/Sample/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4885/SplitProtocol/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4885/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4877/SplitProtocol/Sample/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4877/SplitProtocol/Update/cr
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4877/SplitProtocol/Update/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4877/SplitProtocol/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/$entry
      -- CP-element group 701: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4877/$entry
      -- 
    rr_14033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(701), ack => type_cast_4877_inst_req_0); -- 
    cr_14061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(701), ack => type_cast_4885_inst_req_1); -- 
    rr_14056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(701), ack => type_cast_4885_inst_req_0); -- 
    cr_14038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(701), ack => type_cast_4877_inst_req_1); -- 
    zeropad3D_cp_element_group_701: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_701"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(686) & zeropad3D_CP_2152_elements(688) & zeropad3D_CP_2152_elements(694) & zeropad3D_CP_2152_elements(696) & zeropad3D_CP_2152_elements(698) & zeropad3D_CP_2152_elements(700);
      gj_zeropad3D_cp_element_group_701 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(701), clk => clk, reset => reset); --
    end block;
    -- CP-element group 702:  transition  input  bypass 
    -- CP-element group 702: predecessors 
    -- CP-element group 702: 	1208 
    -- CP-element group 702: successors 
    -- CP-element group 702:  members (3) 
      -- CP-element group 702: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/type_cast_4890_sample_completed_
      -- CP-element group 702: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/type_cast_4890_Sample/ra
      -- CP-element group 702: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/type_cast_4890_Sample/$exit
      -- 
    ra_10181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 702_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4890_inst_ack_0, ack => zeropad3D_CP_2152_elements(702)); -- 
    -- CP-element group 703:  branch  transition  place  input  output  bypass 
    -- CP-element group 703: predecessors 
    -- CP-element group 703: 	1208 
    -- CP-element group 703: successors 
    -- CP-element group 703: 	704 
    -- CP-element group 703: 	705 
    -- CP-element group 703:  members (13) 
      -- CP-element group 703: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898__exit__
      -- CP-element group 703: 	 branch_block_stmt_714/if_stmt_4899__entry__
      -- CP-element group 703: 	 branch_block_stmt_714/R_cmp1567_4900_place
      -- CP-element group 703: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/$exit
      -- CP-element group 703: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/type_cast_4890_Update/ca
      -- CP-element group 703: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/type_cast_4890_update_completed_
      -- CP-element group 703: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/type_cast_4890_Update/$exit
      -- CP-element group 703: 	 branch_block_stmt_714/if_stmt_4899_dead_link/$entry
      -- CP-element group 703: 	 branch_block_stmt_714/if_stmt_4899_eval_test/$entry
      -- CP-element group 703: 	 branch_block_stmt_714/if_stmt_4899_eval_test/$exit
      -- CP-element group 703: 	 branch_block_stmt_714/if_stmt_4899_eval_test/branch_req
      -- CP-element group 703: 	 branch_block_stmt_714/if_stmt_4899_if_link/$entry
      -- CP-element group 703: 	 branch_block_stmt_714/if_stmt_4899_else_link/$entry
      -- 
    ca_10186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 703_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4890_inst_ack_1, ack => zeropad3D_CP_2152_elements(703)); -- 
    branch_req_10194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(703), ack => if_stmt_4899_branch_req_0); -- 
    -- CP-element group 704:  transition  place  input  bypass 
    -- CP-element group 704: predecessors 
    -- CP-element group 704: 	703 
    -- CP-element group 704: successors 
    -- CP-element group 704: 	1209 
    -- CP-element group 704:  members (5) 
      -- CP-element group 704: 	 branch_block_stmt_714/whilex_xbody1562_ifx_xthen1596
      -- CP-element group 704: 	 branch_block_stmt_714/if_stmt_4899_if_link/$exit
      -- CP-element group 704: 	 branch_block_stmt_714/if_stmt_4899_if_link/if_choice_transition
      -- CP-element group 704: 	 branch_block_stmt_714/whilex_xbody1562_ifx_xthen1596_PhiReq/$exit
      -- CP-element group 704: 	 branch_block_stmt_714/whilex_xbody1562_ifx_xthen1596_PhiReq/$entry
      -- 
    if_choice_transition_10199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 704_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4899_branch_ack_1, ack => zeropad3D_CP_2152_elements(704)); -- 
    -- CP-element group 705:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 705: predecessors 
    -- CP-element group 705: 	703 
    -- CP-element group 705: successors 
    -- CP-element group 705: 	706 
    -- CP-element group 705: 	707 
    -- CP-element group 705: 	709 
    -- CP-element group 705:  members (27) 
      -- CP-element group 705: 	 branch_block_stmt_714/merge_stmt_4905__exit__
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924__entry__
      -- CP-element group 705: 	 branch_block_stmt_714/if_stmt_4899_else_link/$exit
      -- CP-element group 705: 	 branch_block_stmt_714/if_stmt_4899_else_link/else_choice_transition
      -- CP-element group 705: 	 branch_block_stmt_714/whilex_xbody1562_lorx_xlhsx_xfalse1569
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/$entry
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_sample_start_
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_update_start_
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_word_address_calculated
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_root_address_calculated
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Sample/$entry
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Sample/word_access_start/$entry
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Sample/word_access_start/word_0/$entry
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Sample/word_access_start/word_0/rr
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Update/$entry
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Update/word_access_complete/$entry
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Update/word_access_complete/word_0/$entry
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Update/word_access_complete/word_0/cr
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/type_cast_4911_update_start_
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/type_cast_4911_Update/$entry
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/type_cast_4911_Update/cr
      -- CP-element group 705: 	 branch_block_stmt_714/whilex_xbody1562_lorx_xlhsx_xfalse1569_PhiReq/$entry
      -- CP-element group 705: 	 branch_block_stmt_714/merge_stmt_4905_PhiReqMerge
      -- CP-element group 705: 	 branch_block_stmt_714/whilex_xbody1562_lorx_xlhsx_xfalse1569_PhiReq/$exit
      -- CP-element group 705: 	 branch_block_stmt_714/merge_stmt_4905_PhiAck/$entry
      -- CP-element group 705: 	 branch_block_stmt_714/merge_stmt_4905_PhiAck/$exit
      -- CP-element group 705: 	 branch_block_stmt_714/merge_stmt_4905_PhiAck/dummy
      -- 
    else_choice_transition_10203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 705_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4899_branch_ack_0, ack => zeropad3D_CP_2152_elements(705)); -- 
    rr_10224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(705), ack => LOAD_row_high_4907_load_0_req_0); -- 
    cr_10235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(705), ack => LOAD_row_high_4907_load_0_req_1); -- 
    cr_10254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(705), ack => type_cast_4911_inst_req_1); -- 
    -- CP-element group 706:  transition  input  bypass 
    -- CP-element group 706: predecessors 
    -- CP-element group 706: 	705 
    -- CP-element group 706: successors 
    -- CP-element group 706:  members (5) 
      -- CP-element group 706: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_sample_completed_
      -- CP-element group 706: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Sample/$exit
      -- CP-element group 706: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Sample/word_access_start/$exit
      -- CP-element group 706: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Sample/word_access_start/word_0/$exit
      -- CP-element group 706: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Sample/word_access_start/word_0/ra
      -- 
    ra_10225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 706_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4907_load_0_ack_0, ack => zeropad3D_CP_2152_elements(706)); -- 
    -- CP-element group 707:  transition  input  output  bypass 
    -- CP-element group 707: predecessors 
    -- CP-element group 707: 	705 
    -- CP-element group 707: successors 
    -- CP-element group 707: 	708 
    -- CP-element group 707:  members (12) 
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_update_completed_
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Update/$exit
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Update/word_access_complete/$exit
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Update/word_access_complete/word_0/$exit
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Update/word_access_complete/word_0/ca
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Update/LOAD_row_high_4907_Merge/$entry
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Update/LOAD_row_high_4907_Merge/$exit
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Update/LOAD_row_high_4907_Merge/merge_req
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/LOAD_row_high_4907_Update/LOAD_row_high_4907_Merge/merge_ack
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/type_cast_4911_sample_start_
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/type_cast_4911_Sample/$entry
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/type_cast_4911_Sample/rr
      -- 
    ca_10236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 707_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4907_load_0_ack_1, ack => zeropad3D_CP_2152_elements(707)); -- 
    rr_10249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(707), ack => type_cast_4911_inst_req_0); -- 
    -- CP-element group 708:  transition  input  bypass 
    -- CP-element group 708: predecessors 
    -- CP-element group 708: 	707 
    -- CP-element group 708: successors 
    -- CP-element group 708:  members (3) 
      -- CP-element group 708: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/type_cast_4911_sample_completed_
      -- CP-element group 708: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/type_cast_4911_Sample/$exit
      -- CP-element group 708: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/type_cast_4911_Sample/ra
      -- 
    ra_10250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 708_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4911_inst_ack_0, ack => zeropad3D_CP_2152_elements(708)); -- 
    -- CP-element group 709:  branch  transition  place  input  output  bypass 
    -- CP-element group 709: predecessors 
    -- CP-element group 709: 	705 
    -- CP-element group 709: successors 
    -- CP-element group 709: 	710 
    -- CP-element group 709: 	711 
    -- CP-element group 709:  members (13) 
      -- CP-element group 709: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924__exit__
      -- CP-element group 709: 	 branch_block_stmt_714/if_stmt_4925__entry__
      -- CP-element group 709: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/$exit
      -- CP-element group 709: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/type_cast_4911_update_completed_
      -- CP-element group 709: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/type_cast_4911_Update/$exit
      -- CP-element group 709: 	 branch_block_stmt_714/assign_stmt_4908_to_assign_stmt_4924/type_cast_4911_Update/ca
      -- CP-element group 709: 	 branch_block_stmt_714/if_stmt_4925_dead_link/$entry
      -- CP-element group 709: 	 branch_block_stmt_714/if_stmt_4925_eval_test/$entry
      -- CP-element group 709: 	 branch_block_stmt_714/if_stmt_4925_eval_test/$exit
      -- CP-element group 709: 	 branch_block_stmt_714/if_stmt_4925_eval_test/branch_req
      -- CP-element group 709: 	 branch_block_stmt_714/R_cmp1577_4926_place
      -- CP-element group 709: 	 branch_block_stmt_714/if_stmt_4925_if_link/$entry
      -- CP-element group 709: 	 branch_block_stmt_714/if_stmt_4925_else_link/$entry
      -- 
    ca_10255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 709_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4911_inst_ack_1, ack => zeropad3D_CP_2152_elements(709)); -- 
    branch_req_10263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(709), ack => if_stmt_4925_branch_req_0); -- 
    -- CP-element group 710:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 710: predecessors 
    -- CP-element group 710: 	709 
    -- CP-element group 710: successors 
    -- CP-element group 710: 	712 
    -- CP-element group 710: 	713 
    -- CP-element group 710:  members (18) 
      -- CP-element group 710: 	 branch_block_stmt_714/merge_stmt_4931__exit__
      -- CP-element group 710: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943__entry__
      -- CP-element group 710: 	 branch_block_stmt_714/if_stmt_4925_if_link/$exit
      -- CP-element group 710: 	 branch_block_stmt_714/if_stmt_4925_if_link/if_choice_transition
      -- CP-element group 710: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1569_lorx_xlhsx_xfalse1579
      -- CP-element group 710: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/$entry
      -- CP-element group 710: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/type_cast_4935_sample_start_
      -- CP-element group 710: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/type_cast_4935_update_start_
      -- CP-element group 710: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/type_cast_4935_Sample/$entry
      -- CP-element group 710: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/type_cast_4935_Sample/rr
      -- CP-element group 710: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/type_cast_4935_Update/$entry
      -- CP-element group 710: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/type_cast_4935_Update/cr
      -- CP-element group 710: 	 branch_block_stmt_714/merge_stmt_4931_PhiReqMerge
      -- CP-element group 710: 	 branch_block_stmt_714/merge_stmt_4931_PhiAck/dummy
      -- CP-element group 710: 	 branch_block_stmt_714/merge_stmt_4931_PhiAck/$exit
      -- CP-element group 710: 	 branch_block_stmt_714/merge_stmt_4931_PhiAck/$entry
      -- CP-element group 710: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1569_lorx_xlhsx_xfalse1579_PhiReq/$exit
      -- CP-element group 710: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1569_lorx_xlhsx_xfalse1579_PhiReq/$entry
      -- 
    if_choice_transition_10268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 710_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4925_branch_ack_1, ack => zeropad3D_CP_2152_elements(710)); -- 
    rr_10285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(710), ack => type_cast_4935_inst_req_0); -- 
    cr_10290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(710), ack => type_cast_4935_inst_req_1); -- 
    -- CP-element group 711:  transition  place  input  bypass 
    -- CP-element group 711: predecessors 
    -- CP-element group 711: 	709 
    -- CP-element group 711: successors 
    -- CP-element group 711: 	1209 
    -- CP-element group 711:  members (5) 
      -- CP-element group 711: 	 branch_block_stmt_714/if_stmt_4925_else_link/$exit
      -- CP-element group 711: 	 branch_block_stmt_714/if_stmt_4925_else_link/else_choice_transition
      -- CP-element group 711: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1569_ifx_xthen1596
      -- CP-element group 711: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1569_ifx_xthen1596_PhiReq/$entry
      -- CP-element group 711: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1569_ifx_xthen1596_PhiReq/$exit
      -- 
    else_choice_transition_10272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 711_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4925_branch_ack_0, ack => zeropad3D_CP_2152_elements(711)); -- 
    -- CP-element group 712:  transition  input  bypass 
    -- CP-element group 712: predecessors 
    -- CP-element group 712: 	710 
    -- CP-element group 712: successors 
    -- CP-element group 712:  members (3) 
      -- CP-element group 712: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/type_cast_4935_sample_completed_
      -- CP-element group 712: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/type_cast_4935_Sample/$exit
      -- CP-element group 712: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/type_cast_4935_Sample/ra
      -- 
    ra_10286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 712_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4935_inst_ack_0, ack => zeropad3D_CP_2152_elements(712)); -- 
    -- CP-element group 713:  branch  transition  place  input  output  bypass 
    -- CP-element group 713: predecessors 
    -- CP-element group 713: 	710 
    -- CP-element group 713: successors 
    -- CP-element group 713: 	714 
    -- CP-element group 713: 	715 
    -- CP-element group 713:  members (13) 
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943__exit__
      -- CP-element group 713: 	 branch_block_stmt_714/if_stmt_4944__entry__
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/$exit
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/type_cast_4935_update_completed_
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/type_cast_4935_Update/$exit
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4936_to_assign_stmt_4943/type_cast_4935_Update/ca
      -- CP-element group 713: 	 branch_block_stmt_714/if_stmt_4944_dead_link/$entry
      -- CP-element group 713: 	 branch_block_stmt_714/if_stmt_4944_eval_test/$entry
      -- CP-element group 713: 	 branch_block_stmt_714/if_stmt_4944_eval_test/$exit
      -- CP-element group 713: 	 branch_block_stmt_714/if_stmt_4944_eval_test/branch_req
      -- CP-element group 713: 	 branch_block_stmt_714/R_cmp1584_4945_place
      -- CP-element group 713: 	 branch_block_stmt_714/if_stmt_4944_if_link/$entry
      -- CP-element group 713: 	 branch_block_stmt_714/if_stmt_4944_else_link/$entry
      -- 
    ca_10291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 713_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4935_inst_ack_1, ack => zeropad3D_CP_2152_elements(713)); -- 
    branch_req_10299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(713), ack => if_stmt_4944_branch_req_0); -- 
    -- CP-element group 714:  transition  place  input  bypass 
    -- CP-element group 714: predecessors 
    -- CP-element group 714: 	713 
    -- CP-element group 714: successors 
    -- CP-element group 714: 	1209 
    -- CP-element group 714:  members (5) 
      -- CP-element group 714: 	 branch_block_stmt_714/if_stmt_4944_if_link/$exit
      -- CP-element group 714: 	 branch_block_stmt_714/if_stmt_4944_if_link/if_choice_transition
      -- CP-element group 714: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1579_ifx_xthen1596
      -- CP-element group 714: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1579_ifx_xthen1596_PhiReq/$exit
      -- CP-element group 714: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1579_ifx_xthen1596_PhiReq/$entry
      -- 
    if_choice_transition_10304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 714_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4944_branch_ack_1, ack => zeropad3D_CP_2152_elements(714)); -- 
    -- CP-element group 715:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 715: predecessors 
    -- CP-element group 715: 	713 
    -- CP-element group 715: successors 
    -- CP-element group 715: 	716 
    -- CP-element group 715: 	717 
    -- CP-element group 715: 	719 
    -- CP-element group 715:  members (27) 
      -- CP-element group 715: 	 branch_block_stmt_714/merge_stmt_4950__exit__
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969__entry__
      -- CP-element group 715: 	 branch_block_stmt_714/if_stmt_4944_else_link/$exit
      -- CP-element group 715: 	 branch_block_stmt_714/if_stmt_4944_else_link/else_choice_transition
      -- CP-element group 715: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1579_lorx_xlhsx_xfalse1586
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/$entry
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_sample_start_
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_update_start_
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_word_address_calculated
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_root_address_calculated
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Sample/$entry
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Sample/word_access_start/$entry
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Sample/word_access_start/word_0/$entry
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Sample/word_access_start/word_0/rr
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Update/$entry
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Update/word_access_complete/$entry
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Update/word_access_complete/word_0/$entry
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Update/word_access_complete/word_0/cr
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/type_cast_4956_update_start_
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/type_cast_4956_Update/$entry
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/type_cast_4956_Update/cr
      -- CP-element group 715: 	 branch_block_stmt_714/merge_stmt_4950_PhiReqMerge
      -- CP-element group 715: 	 branch_block_stmt_714/merge_stmt_4950_PhiAck/dummy
      -- CP-element group 715: 	 branch_block_stmt_714/merge_stmt_4950_PhiAck/$exit
      -- CP-element group 715: 	 branch_block_stmt_714/merge_stmt_4950_PhiAck/$entry
      -- CP-element group 715: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1579_lorx_xlhsx_xfalse1586_PhiReq/$exit
      -- CP-element group 715: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1579_lorx_xlhsx_xfalse1586_PhiReq/$entry
      -- 
    else_choice_transition_10308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 715_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4944_branch_ack_0, ack => zeropad3D_CP_2152_elements(715)); -- 
    rr_10329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(715), ack => LOAD_col_high_4952_load_0_req_0); -- 
    cr_10340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(715), ack => LOAD_col_high_4952_load_0_req_1); -- 
    cr_10359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(715), ack => type_cast_4956_inst_req_1); -- 
    -- CP-element group 716:  transition  input  bypass 
    -- CP-element group 716: predecessors 
    -- CP-element group 716: 	715 
    -- CP-element group 716: successors 
    -- CP-element group 716:  members (5) 
      -- CP-element group 716: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_sample_completed_
      -- CP-element group 716: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Sample/$exit
      -- CP-element group 716: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Sample/word_access_start/$exit
      -- CP-element group 716: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Sample/word_access_start/word_0/$exit
      -- CP-element group 716: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Sample/word_access_start/word_0/ra
      -- 
    ra_10330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 716_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4952_load_0_ack_0, ack => zeropad3D_CP_2152_elements(716)); -- 
    -- CP-element group 717:  transition  input  output  bypass 
    -- CP-element group 717: predecessors 
    -- CP-element group 717: 	715 
    -- CP-element group 717: successors 
    -- CP-element group 717: 	718 
    -- CP-element group 717:  members (12) 
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_update_completed_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Update/$exit
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Update/word_access_complete/$exit
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Update/word_access_complete/word_0/$exit
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Update/word_access_complete/word_0/ca
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Update/LOAD_col_high_4952_Merge/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Update/LOAD_col_high_4952_Merge/$exit
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Update/LOAD_col_high_4952_Merge/merge_req
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/LOAD_col_high_4952_Update/LOAD_col_high_4952_Merge/merge_ack
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/type_cast_4956_sample_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/type_cast_4956_Sample/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/type_cast_4956_Sample/rr
      -- 
    ca_10341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 717_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4952_load_0_ack_1, ack => zeropad3D_CP_2152_elements(717)); -- 
    rr_10354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => type_cast_4956_inst_req_0); -- 
    -- CP-element group 718:  transition  input  bypass 
    -- CP-element group 718: predecessors 
    -- CP-element group 718: 	717 
    -- CP-element group 718: successors 
    -- CP-element group 718:  members (3) 
      -- CP-element group 718: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/type_cast_4956_sample_completed_
      -- CP-element group 718: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/type_cast_4956_Sample/$exit
      -- CP-element group 718: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/type_cast_4956_Sample/ra
      -- 
    ra_10355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 718_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4956_inst_ack_0, ack => zeropad3D_CP_2152_elements(718)); -- 
    -- CP-element group 719:  branch  transition  place  input  output  bypass 
    -- CP-element group 719: predecessors 
    -- CP-element group 719: 	715 
    -- CP-element group 719: successors 
    -- CP-element group 719: 	720 
    -- CP-element group 719: 	721 
    -- CP-element group 719:  members (13) 
      -- CP-element group 719: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969__exit__
      -- CP-element group 719: 	 branch_block_stmt_714/if_stmt_4970__entry__
      -- CP-element group 719: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/$exit
      -- CP-element group 719: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/type_cast_4956_update_completed_
      -- CP-element group 719: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/type_cast_4956_Update/$exit
      -- CP-element group 719: 	 branch_block_stmt_714/assign_stmt_4953_to_assign_stmt_4969/type_cast_4956_Update/ca
      -- CP-element group 719: 	 branch_block_stmt_714/if_stmt_4970_dead_link/$entry
      -- CP-element group 719: 	 branch_block_stmt_714/if_stmt_4970_eval_test/$entry
      -- CP-element group 719: 	 branch_block_stmt_714/if_stmt_4970_eval_test/$exit
      -- CP-element group 719: 	 branch_block_stmt_714/if_stmt_4970_eval_test/branch_req
      -- CP-element group 719: 	 branch_block_stmt_714/R_cmp1594_4971_place
      -- CP-element group 719: 	 branch_block_stmt_714/if_stmt_4970_if_link/$entry
      -- CP-element group 719: 	 branch_block_stmt_714/if_stmt_4970_else_link/$entry
      -- 
    ca_10360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 719_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4956_inst_ack_1, ack => zeropad3D_CP_2152_elements(719)); -- 
    branch_req_10368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(719), ack => if_stmt_4970_branch_req_0); -- 
    -- CP-element group 720:  fork  transition  place  input  output  bypass 
    -- CP-element group 720: predecessors 
    -- CP-element group 720: 	719 
    -- CP-element group 720: successors 
    -- CP-element group 720: 	736 
    -- CP-element group 720: 	737 
    -- CP-element group 720: 	739 
    -- CP-element group 720: 	741 
    -- CP-element group 720: 	743 
    -- CP-element group 720: 	745 
    -- CP-element group 720: 	747 
    -- CP-element group 720: 	749 
    -- CP-element group 720: 	751 
    -- CP-element group 720: 	754 
    -- CP-element group 720:  members (46) 
      -- CP-element group 720: 	 branch_block_stmt_714/merge_stmt_5034__exit__
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139__entry__
      -- CP-element group 720: 	 branch_block_stmt_714/if_stmt_4970_if_link/$exit
      -- CP-element group 720: 	 branch_block_stmt_714/if_stmt_4970_if_link/if_choice_transition
      -- CP-element group 720: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1586_ifx_xelse1617
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5038_sample_start_
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5038_update_start_
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5038_Sample/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5038_Sample/rr
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5038_Update/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5038_Update/cr
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5102_update_start_
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5102_Update/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5102_Update/cr
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5109_update_start_
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_final_index_sum_regn_update_start
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_final_index_sum_regn_Update/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_final_index_sum_regn_Update/req
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5109_complete/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5109_complete/req
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_update_start_
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Update/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Update/word_access_complete/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Update/word_access_complete/word_0/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Update/word_access_complete/word_0/cr
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5127_update_start_
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5127_Update/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5127_Update/cr
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5134_update_start_
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_final_index_sum_regn_update_start
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_final_index_sum_regn_Update/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_final_index_sum_regn_Update/req
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5134_complete/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5134_complete/req
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_update_start_
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Update/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Update/word_access_complete/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Update/word_access_complete/word_0/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Update/word_access_complete/word_0/cr
      -- CP-element group 720: 	 branch_block_stmt_714/merge_stmt_5034_PhiReqMerge
      -- CP-element group 720: 	 branch_block_stmt_714/merge_stmt_5034_PhiAck/dummy
      -- CP-element group 720: 	 branch_block_stmt_714/merge_stmt_5034_PhiAck/$exit
      -- CP-element group 720: 	 branch_block_stmt_714/merge_stmt_5034_PhiAck/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1586_ifx_xelse1617_PhiReq/$exit
      -- CP-element group 720: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1586_ifx_xelse1617_PhiReq/$entry
      -- 
    if_choice_transition_10373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 720_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4970_branch_ack_1, ack => zeropad3D_CP_2152_elements(720)); -- 
    rr_10531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(720), ack => type_cast_5038_inst_req_0); -- 
    cr_10536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(720), ack => type_cast_5038_inst_req_1); -- 
    cr_10550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(720), ack => type_cast_5102_inst_req_1); -- 
    req_10581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(720), ack => array_obj_ref_5108_index_offset_req_1); -- 
    req_10596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(720), ack => addr_of_5109_final_reg_req_1); -- 
    cr_10641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(720), ack => ptr_deref_5113_load_0_req_1); -- 
    cr_10660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(720), ack => type_cast_5127_inst_req_1); -- 
    req_10691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(720), ack => array_obj_ref_5133_index_offset_req_1); -- 
    req_10706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(720), ack => addr_of_5134_final_reg_req_1); -- 
    cr_10756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(720), ack => ptr_deref_5137_store_0_req_1); -- 
    -- CP-element group 721:  transition  place  input  bypass 
    -- CP-element group 721: predecessors 
    -- CP-element group 721: 	719 
    -- CP-element group 721: successors 
    -- CP-element group 721: 	1209 
    -- CP-element group 721:  members (5) 
      -- CP-element group 721: 	 branch_block_stmt_714/if_stmt_4970_else_link/$exit
      -- CP-element group 721: 	 branch_block_stmt_714/if_stmt_4970_else_link/else_choice_transition
      -- CP-element group 721: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1586_ifx_xthen1596
      -- CP-element group 721: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1586_ifx_xthen1596_PhiReq/$exit
      -- CP-element group 721: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1586_ifx_xthen1596_PhiReq/$entry
      -- 
    else_choice_transition_10377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 721_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4970_branch_ack_0, ack => zeropad3D_CP_2152_elements(721)); -- 
    -- CP-element group 722:  transition  input  bypass 
    -- CP-element group 722: predecessors 
    -- CP-element group 722: 	1209 
    -- CP-element group 722: successors 
    -- CP-element group 722:  members (3) 
      -- CP-element group 722: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4980_sample_completed_
      -- CP-element group 722: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4980_Sample/$exit
      -- CP-element group 722: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4980_Sample/ra
      -- 
    ra_10391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 722_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4980_inst_ack_0, ack => zeropad3D_CP_2152_elements(722)); -- 
    -- CP-element group 723:  transition  input  bypass 
    -- CP-element group 723: predecessors 
    -- CP-element group 723: 	1209 
    -- CP-element group 723: successors 
    -- CP-element group 723: 	726 
    -- CP-element group 723:  members (3) 
      -- CP-element group 723: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4980_update_completed_
      -- CP-element group 723: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4980_Update/$exit
      -- CP-element group 723: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4980_Update/ca
      -- 
    ca_10396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 723_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4980_inst_ack_1, ack => zeropad3D_CP_2152_elements(723)); -- 
    -- CP-element group 724:  transition  input  bypass 
    -- CP-element group 724: predecessors 
    -- CP-element group 724: 	1209 
    -- CP-element group 724: successors 
    -- CP-element group 724:  members (3) 
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4985_sample_completed_
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4985_Sample/$exit
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4985_Sample/ra
      -- 
    ra_10405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 724_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4985_inst_ack_0, ack => zeropad3D_CP_2152_elements(724)); -- 
    -- CP-element group 725:  transition  input  bypass 
    -- CP-element group 725: predecessors 
    -- CP-element group 725: 	1209 
    -- CP-element group 725: successors 
    -- CP-element group 725: 	726 
    -- CP-element group 725:  members (3) 
      -- CP-element group 725: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4985_update_completed_
      -- CP-element group 725: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4985_Update/$exit
      -- CP-element group 725: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4985_Update/ca
      -- 
    ca_10410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 725_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4985_inst_ack_1, ack => zeropad3D_CP_2152_elements(725)); -- 
    -- CP-element group 726:  join  transition  output  bypass 
    -- CP-element group 726: predecessors 
    -- CP-element group 726: 	723 
    -- CP-element group 726: 	725 
    -- CP-element group 726: successors 
    -- CP-element group 726: 	727 
    -- CP-element group 726:  members (3) 
      -- CP-element group 726: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_5019_sample_start_
      -- CP-element group 726: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_5019_Sample/$entry
      -- CP-element group 726: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_5019_Sample/rr
      -- 
    rr_10418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(726), ack => type_cast_5019_inst_req_0); -- 
    zeropad3D_cp_element_group_726: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_726"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(723) & zeropad3D_CP_2152_elements(725);
      gj_zeropad3D_cp_element_group_726 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(726), clk => clk, reset => reset); --
    end block;
    -- CP-element group 727:  transition  input  bypass 
    -- CP-element group 727: predecessors 
    -- CP-element group 727: 	726 
    -- CP-element group 727: successors 
    -- CP-element group 727:  members (3) 
      -- CP-element group 727: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_5019_sample_completed_
      -- CP-element group 727: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_5019_Sample/$exit
      -- CP-element group 727: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_5019_Sample/ra
      -- 
    ra_10419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 727_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5019_inst_ack_0, ack => zeropad3D_CP_2152_elements(727)); -- 
    -- CP-element group 728:  transition  input  output  bypass 
    -- CP-element group 728: predecessors 
    -- CP-element group 728: 	1209 
    -- CP-element group 728: successors 
    -- CP-element group 728: 	729 
    -- CP-element group 728:  members (16) 
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_5019_update_completed_
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_5019_Update/$exit
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_5019_Update/ca
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_index_resized_1
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_index_scaled_1
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_index_computed_1
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_index_resize_1/$entry
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_index_resize_1/$exit
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_index_resize_1/index_resize_req
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_index_resize_1/index_resize_ack
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_index_scale_1/$entry
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_index_scale_1/$exit
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_index_scale_1/scale_rename_req
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_index_scale_1/scale_rename_ack
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_final_index_sum_regn_Sample/$entry
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_final_index_sum_regn_Sample/req
      -- 
    ca_10424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 728_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5019_inst_ack_1, ack => zeropad3D_CP_2152_elements(728)); -- 
    req_10449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(728), ack => array_obj_ref_5025_index_offset_req_0); -- 
    -- CP-element group 729:  transition  input  bypass 
    -- CP-element group 729: predecessors 
    -- CP-element group 729: 	728 
    -- CP-element group 729: successors 
    -- CP-element group 729: 	735 
    -- CP-element group 729:  members (3) 
      -- CP-element group 729: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_final_index_sum_regn_sample_complete
      -- CP-element group 729: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_final_index_sum_regn_Sample/$exit
      -- CP-element group 729: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_final_index_sum_regn_Sample/ack
      -- 
    ack_10450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 729_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_5025_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(729)); -- 
    -- CP-element group 730:  transition  input  output  bypass 
    -- CP-element group 730: predecessors 
    -- CP-element group 730: 	1209 
    -- CP-element group 730: successors 
    -- CP-element group 730: 	731 
    -- CP-element group 730:  members (11) 
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/addr_of_5026_sample_start_
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_root_address_calculated
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_offset_calculated
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_final_index_sum_regn_Update/$exit
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_final_index_sum_regn_Update/ack
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_base_plus_offset/$entry
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_base_plus_offset/$exit
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_base_plus_offset/sum_rename_req
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_base_plus_offset/sum_rename_ack
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/addr_of_5026_request/$entry
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/addr_of_5026_request/req
      -- 
    ack_10455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 730_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_5025_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(730)); -- 
    req_10464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(730), ack => addr_of_5026_final_reg_req_0); -- 
    -- CP-element group 731:  transition  input  bypass 
    -- CP-element group 731: predecessors 
    -- CP-element group 731: 	730 
    -- CP-element group 731: successors 
    -- CP-element group 731:  members (3) 
      -- CP-element group 731: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/addr_of_5026_sample_completed_
      -- CP-element group 731: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/addr_of_5026_request/$exit
      -- CP-element group 731: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/addr_of_5026_request/ack
      -- 
    ack_10465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 731_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_5026_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(731)); -- 
    -- CP-element group 732:  join  fork  transition  input  output  bypass 
    -- CP-element group 732: predecessors 
    -- CP-element group 732: 	1209 
    -- CP-element group 732: successors 
    -- CP-element group 732: 	733 
    -- CP-element group 732:  members (28) 
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/addr_of_5026_update_completed_
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/addr_of_5026_complete/$exit
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/addr_of_5026_complete/ack
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_sample_start_
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_base_address_calculated
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_word_address_calculated
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_root_address_calculated
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_base_address_resized
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_base_addr_resize/$entry
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_base_addr_resize/$exit
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_base_addr_resize/base_resize_req
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_base_addr_resize/base_resize_ack
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_base_plus_offset/$entry
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_base_plus_offset/$exit
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_base_plus_offset/sum_rename_req
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_base_plus_offset/sum_rename_ack
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_word_addrgen/$entry
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_word_addrgen/$exit
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_word_addrgen/root_register_req
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_word_addrgen/root_register_ack
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Sample/$entry
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Sample/ptr_deref_5029_Split/$entry
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Sample/ptr_deref_5029_Split/$exit
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Sample/ptr_deref_5029_Split/split_req
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Sample/ptr_deref_5029_Split/split_ack
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Sample/word_access_start/$entry
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Sample/word_access_start/word_0/$entry
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Sample/word_access_start/word_0/rr
      -- 
    ack_10470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 732_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_5026_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(732)); -- 
    rr_10508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(732), ack => ptr_deref_5029_store_0_req_0); -- 
    -- CP-element group 733:  transition  input  bypass 
    -- CP-element group 733: predecessors 
    -- CP-element group 733: 	732 
    -- CP-element group 733: successors 
    -- CP-element group 733:  members (5) 
      -- CP-element group 733: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_sample_completed_
      -- CP-element group 733: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Sample/$exit
      -- CP-element group 733: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Sample/word_access_start/$exit
      -- CP-element group 733: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Sample/word_access_start/word_0/$exit
      -- CP-element group 733: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Sample/word_access_start/word_0/ra
      -- 
    ra_10509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 733_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_5029_store_0_ack_0, ack => zeropad3D_CP_2152_elements(733)); -- 
    -- CP-element group 734:  transition  input  bypass 
    -- CP-element group 734: predecessors 
    -- CP-element group 734: 	1209 
    -- CP-element group 734: successors 
    -- CP-element group 734: 	735 
    -- CP-element group 734:  members (5) 
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_update_completed_
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Update/$exit
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Update/word_access_complete/$exit
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Update/word_access_complete/word_0/$exit
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Update/word_access_complete/word_0/ca
      -- 
    ca_10520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 734_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_5029_store_0_ack_1, ack => zeropad3D_CP_2152_elements(734)); -- 
    -- CP-element group 735:  join  transition  place  bypass 
    -- CP-element group 735: predecessors 
    -- CP-element group 735: 	729 
    -- CP-element group 735: 	734 
    -- CP-element group 735: successors 
    -- CP-element group 735: 	1210 
    -- CP-element group 735:  members (5) 
      -- CP-element group 735: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032__exit__
      -- CP-element group 735: 	 branch_block_stmt_714/ifx_xthen1596_ifx_xend1665
      -- CP-element group 735: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/$exit
      -- CP-element group 735: 	 branch_block_stmt_714/ifx_xthen1596_ifx_xend1665_PhiReq/$exit
      -- CP-element group 735: 	 branch_block_stmt_714/ifx_xthen1596_ifx_xend1665_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_735: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_735"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(729) & zeropad3D_CP_2152_elements(734);
      gj_zeropad3D_cp_element_group_735 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(735), clk => clk, reset => reset); --
    end block;
    -- CP-element group 736:  transition  input  bypass 
    -- CP-element group 736: predecessors 
    -- CP-element group 736: 	720 
    -- CP-element group 736: successors 
    -- CP-element group 736:  members (3) 
      -- CP-element group 736: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5038_sample_completed_
      -- CP-element group 736: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5038_Sample/$exit
      -- CP-element group 736: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5038_Sample/ra
      -- 
    ra_10532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 736_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5038_inst_ack_0, ack => zeropad3D_CP_2152_elements(736)); -- 
    -- CP-element group 737:  fork  transition  input  output  bypass 
    -- CP-element group 737: predecessors 
    -- CP-element group 737: 	720 
    -- CP-element group 737: successors 
    -- CP-element group 737: 	738 
    -- CP-element group 737: 	746 
    -- CP-element group 737:  members (9) 
      -- CP-element group 737: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5038_update_completed_
      -- CP-element group 737: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5038_Update/$exit
      -- CP-element group 737: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5038_Update/ca
      -- CP-element group 737: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5102_sample_start_
      -- CP-element group 737: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5102_Sample/$entry
      -- CP-element group 737: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5102_Sample/rr
      -- CP-element group 737: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5127_sample_start_
      -- CP-element group 737: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5127_Sample/$entry
      -- CP-element group 737: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5127_Sample/rr
      -- 
    ca_10537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 737_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5038_inst_ack_1, ack => zeropad3D_CP_2152_elements(737)); -- 
    rr_10545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(737), ack => type_cast_5102_inst_req_0); -- 
    rr_10655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(737), ack => type_cast_5127_inst_req_0); -- 
    -- CP-element group 738:  transition  input  bypass 
    -- CP-element group 738: predecessors 
    -- CP-element group 738: 	737 
    -- CP-element group 738: successors 
    -- CP-element group 738:  members (3) 
      -- CP-element group 738: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5102_sample_completed_
      -- CP-element group 738: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5102_Sample/$exit
      -- CP-element group 738: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5102_Sample/ra
      -- 
    ra_10546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 738_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5102_inst_ack_0, ack => zeropad3D_CP_2152_elements(738)); -- 
    -- CP-element group 739:  transition  input  output  bypass 
    -- CP-element group 739: predecessors 
    -- CP-element group 739: 	720 
    -- CP-element group 739: successors 
    -- CP-element group 739: 	740 
    -- CP-element group 739:  members (16) 
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5102_update_completed_
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5102_Update/$exit
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5102_Update/ca
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_index_resized_1
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_index_scaled_1
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_index_computed_1
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_index_resize_1/$entry
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_index_resize_1/$exit
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_index_resize_1/index_resize_req
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_index_resize_1/index_resize_ack
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_index_scale_1/$entry
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_index_scale_1/$exit
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_index_scale_1/scale_rename_req
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_index_scale_1/scale_rename_ack
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_final_index_sum_regn_Sample/$entry
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_final_index_sum_regn_Sample/req
      -- 
    ca_10551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 739_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5102_inst_ack_1, ack => zeropad3D_CP_2152_elements(739)); -- 
    req_10576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(739), ack => array_obj_ref_5108_index_offset_req_0); -- 
    -- CP-element group 740:  transition  input  bypass 
    -- CP-element group 740: predecessors 
    -- CP-element group 740: 	739 
    -- CP-element group 740: successors 
    -- CP-element group 740: 	755 
    -- CP-element group 740:  members (3) 
      -- CP-element group 740: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_final_index_sum_regn_sample_complete
      -- CP-element group 740: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_final_index_sum_regn_Sample/$exit
      -- CP-element group 740: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_final_index_sum_regn_Sample/ack
      -- 
    ack_10577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 740_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_5108_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(740)); -- 
    -- CP-element group 741:  transition  input  output  bypass 
    -- CP-element group 741: predecessors 
    -- CP-element group 741: 	720 
    -- CP-element group 741: successors 
    -- CP-element group 741: 	742 
    -- CP-element group 741:  members (11) 
      -- CP-element group 741: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5109_sample_start_
      -- CP-element group 741: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_root_address_calculated
      -- CP-element group 741: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_offset_calculated
      -- CP-element group 741: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_final_index_sum_regn_Update/$exit
      -- CP-element group 741: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_final_index_sum_regn_Update/ack
      -- CP-element group 741: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_base_plus_offset/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_base_plus_offset/$exit
      -- CP-element group 741: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_base_plus_offset/sum_rename_req
      -- CP-element group 741: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5108_base_plus_offset/sum_rename_ack
      -- CP-element group 741: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5109_request/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5109_request/req
      -- 
    ack_10582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 741_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_5108_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(741)); -- 
    req_10591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(741), ack => addr_of_5109_final_reg_req_0); -- 
    -- CP-element group 742:  transition  input  bypass 
    -- CP-element group 742: predecessors 
    -- CP-element group 742: 	741 
    -- CP-element group 742: successors 
    -- CP-element group 742:  members (3) 
      -- CP-element group 742: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5109_sample_completed_
      -- CP-element group 742: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5109_request/$exit
      -- CP-element group 742: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5109_request/ack
      -- 
    ack_10592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 742_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_5109_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(742)); -- 
    -- CP-element group 743:  join  fork  transition  input  output  bypass 
    -- CP-element group 743: predecessors 
    -- CP-element group 743: 	720 
    -- CP-element group 743: successors 
    -- CP-element group 743: 	744 
    -- CP-element group 743:  members (24) 
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5109_update_completed_
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5109_complete/$exit
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5109_complete/ack
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_sample_start_
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_base_address_calculated
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_word_address_calculated
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_root_address_calculated
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_base_address_resized
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_base_addr_resize/$entry
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_base_addr_resize/$exit
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_base_addr_resize/base_resize_req
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_base_addr_resize/base_resize_ack
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_base_plus_offset/$entry
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_base_plus_offset/$exit
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_base_plus_offset/sum_rename_req
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_base_plus_offset/sum_rename_ack
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_word_addrgen/$entry
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_word_addrgen/$exit
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_word_addrgen/root_register_req
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_word_addrgen/root_register_ack
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Sample/$entry
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Sample/word_access_start/$entry
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Sample/word_access_start/word_0/$entry
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Sample/word_access_start/word_0/rr
      -- 
    ack_10597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 743_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_5109_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(743)); -- 
    rr_10630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(743), ack => ptr_deref_5113_load_0_req_0); -- 
    -- CP-element group 744:  transition  input  bypass 
    -- CP-element group 744: predecessors 
    -- CP-element group 744: 	743 
    -- CP-element group 744: successors 
    -- CP-element group 744:  members (5) 
      -- CP-element group 744: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_sample_completed_
      -- CP-element group 744: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Sample/$exit
      -- CP-element group 744: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Sample/word_access_start/$exit
      -- CP-element group 744: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Sample/word_access_start/word_0/$exit
      -- CP-element group 744: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Sample/word_access_start/word_0/ra
      -- 
    ra_10631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 744_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_5113_load_0_ack_0, ack => zeropad3D_CP_2152_elements(744)); -- 
    -- CP-element group 745:  transition  input  bypass 
    -- CP-element group 745: predecessors 
    -- CP-element group 745: 	720 
    -- CP-element group 745: successors 
    -- CP-element group 745: 	752 
    -- CP-element group 745:  members (9) 
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_update_completed_
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Update/$exit
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Update/word_access_complete/$exit
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Update/word_access_complete/word_0/$exit
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Update/word_access_complete/word_0/ca
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Update/ptr_deref_5113_Merge/$entry
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Update/ptr_deref_5113_Merge/$exit
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Update/ptr_deref_5113_Merge/merge_req
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5113_Update/ptr_deref_5113_Merge/merge_ack
      -- 
    ca_10642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 745_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_5113_load_0_ack_1, ack => zeropad3D_CP_2152_elements(745)); -- 
    -- CP-element group 746:  transition  input  bypass 
    -- CP-element group 746: predecessors 
    -- CP-element group 746: 	737 
    -- CP-element group 746: successors 
    -- CP-element group 746:  members (3) 
      -- CP-element group 746: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5127_sample_completed_
      -- CP-element group 746: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5127_Sample/$exit
      -- CP-element group 746: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5127_Sample/ra
      -- 
    ra_10656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 746_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5127_inst_ack_0, ack => zeropad3D_CP_2152_elements(746)); -- 
    -- CP-element group 747:  transition  input  output  bypass 
    -- CP-element group 747: predecessors 
    -- CP-element group 747: 	720 
    -- CP-element group 747: successors 
    -- CP-element group 747: 	748 
    -- CP-element group 747:  members (16) 
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5127_update_completed_
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5127_Update/$exit
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/type_cast_5127_Update/ca
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_index_resized_1
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_index_scaled_1
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_index_computed_1
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_index_resize_1/$entry
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_index_resize_1/$exit
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_index_resize_1/index_resize_req
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_index_resize_1/index_resize_ack
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_index_scale_1/$entry
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_index_scale_1/$exit
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_index_scale_1/scale_rename_req
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_index_scale_1/scale_rename_ack
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_final_index_sum_regn_Sample/$entry
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_final_index_sum_regn_Sample/req
      -- 
    ca_10661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 747_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5127_inst_ack_1, ack => zeropad3D_CP_2152_elements(747)); -- 
    req_10686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(747), ack => array_obj_ref_5133_index_offset_req_0); -- 
    -- CP-element group 748:  transition  input  bypass 
    -- CP-element group 748: predecessors 
    -- CP-element group 748: 	747 
    -- CP-element group 748: successors 
    -- CP-element group 748: 	755 
    -- CP-element group 748:  members (3) 
      -- CP-element group 748: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_final_index_sum_regn_sample_complete
      -- CP-element group 748: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_final_index_sum_regn_Sample/$exit
      -- CP-element group 748: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_final_index_sum_regn_Sample/ack
      -- 
    ack_10687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 748_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_5133_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(748)); -- 
    -- CP-element group 749:  transition  input  output  bypass 
    -- CP-element group 749: predecessors 
    -- CP-element group 749: 	720 
    -- CP-element group 749: successors 
    -- CP-element group 749: 	750 
    -- CP-element group 749:  members (11) 
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5134_sample_start_
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_root_address_calculated
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_offset_calculated
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_final_index_sum_regn_Update/$exit
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_final_index_sum_regn_Update/ack
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_base_plus_offset/$entry
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_base_plus_offset/$exit
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_base_plus_offset/sum_rename_req
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/array_obj_ref_5133_base_plus_offset/sum_rename_ack
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5134_request/$entry
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5134_request/req
      -- 
    ack_10692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 749_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_5133_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(749)); -- 
    req_10701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(749), ack => addr_of_5134_final_reg_req_0); -- 
    -- CP-element group 750:  transition  input  bypass 
    -- CP-element group 750: predecessors 
    -- CP-element group 750: 	749 
    -- CP-element group 750: successors 
    -- CP-element group 750:  members (3) 
      -- CP-element group 750: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5134_sample_completed_
      -- CP-element group 750: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5134_request/$exit
      -- CP-element group 750: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5134_request/ack
      -- 
    ack_10702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 750_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_5134_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(750)); -- 
    -- CP-element group 751:  fork  transition  input  bypass 
    -- CP-element group 751: predecessors 
    -- CP-element group 751: 	720 
    -- CP-element group 751: successors 
    -- CP-element group 751: 	752 
    -- CP-element group 751:  members (19) 
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5134_update_completed_
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5134_complete/$exit
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/addr_of_5134_complete/ack
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_base_address_calculated
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_word_address_calculated
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_root_address_calculated
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_base_address_resized
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_base_addr_resize/$entry
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_base_addr_resize/$exit
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_base_addr_resize/base_resize_req
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_base_addr_resize/base_resize_ack
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_base_plus_offset/$entry
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_base_plus_offset/$exit
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_base_plus_offset/sum_rename_req
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_base_plus_offset/sum_rename_ack
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_word_addrgen/$entry
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_word_addrgen/$exit
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_word_addrgen/root_register_req
      -- CP-element group 751: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_word_addrgen/root_register_ack
      -- 
    ack_10707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 751_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_5134_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(751)); -- 
    -- CP-element group 752:  join  transition  output  bypass 
    -- CP-element group 752: predecessors 
    -- CP-element group 752: 	745 
    -- CP-element group 752: 	751 
    -- CP-element group 752: successors 
    -- CP-element group 752: 	753 
    -- CP-element group 752:  members (9) 
      -- CP-element group 752: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_sample_start_
      -- CP-element group 752: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Sample/$entry
      -- CP-element group 752: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Sample/ptr_deref_5137_Split/$entry
      -- CP-element group 752: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Sample/ptr_deref_5137_Split/$exit
      -- CP-element group 752: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Sample/ptr_deref_5137_Split/split_req
      -- CP-element group 752: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Sample/ptr_deref_5137_Split/split_ack
      -- CP-element group 752: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Sample/word_access_start/$entry
      -- CP-element group 752: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Sample/word_access_start/word_0/$entry
      -- CP-element group 752: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Sample/word_access_start/word_0/rr
      -- 
    rr_10745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(752), ack => ptr_deref_5137_store_0_req_0); -- 
    zeropad3D_cp_element_group_752: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_752"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(745) & zeropad3D_CP_2152_elements(751);
      gj_zeropad3D_cp_element_group_752 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(752), clk => clk, reset => reset); --
    end block;
    -- CP-element group 753:  transition  input  bypass 
    -- CP-element group 753: predecessors 
    -- CP-element group 753: 	752 
    -- CP-element group 753: successors 
    -- CP-element group 753:  members (5) 
      -- CP-element group 753: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_sample_completed_
      -- CP-element group 753: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Sample/$exit
      -- CP-element group 753: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Sample/word_access_start/$exit
      -- CP-element group 753: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Sample/word_access_start/word_0/$exit
      -- CP-element group 753: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Sample/word_access_start/word_0/ra
      -- 
    ra_10746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 753_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_5137_store_0_ack_0, ack => zeropad3D_CP_2152_elements(753)); -- 
    -- CP-element group 754:  transition  input  bypass 
    -- CP-element group 754: predecessors 
    -- CP-element group 754: 	720 
    -- CP-element group 754: successors 
    -- CP-element group 754: 	755 
    -- CP-element group 754:  members (5) 
      -- CP-element group 754: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_update_completed_
      -- CP-element group 754: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Update/$exit
      -- CP-element group 754: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Update/word_access_complete/$exit
      -- CP-element group 754: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Update/word_access_complete/word_0/$exit
      -- CP-element group 754: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/ptr_deref_5137_Update/word_access_complete/word_0/ca
      -- 
    ca_10757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 754_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_5137_store_0_ack_1, ack => zeropad3D_CP_2152_elements(754)); -- 
    -- CP-element group 755:  join  transition  place  bypass 
    -- CP-element group 755: predecessors 
    -- CP-element group 755: 	740 
    -- CP-element group 755: 	748 
    -- CP-element group 755: 	754 
    -- CP-element group 755: successors 
    -- CP-element group 755: 	1210 
    -- CP-element group 755:  members (5) 
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139__exit__
      -- CP-element group 755: 	 branch_block_stmt_714/ifx_xelse1617_ifx_xend1665
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_5039_to_assign_stmt_5139/$exit
      -- CP-element group 755: 	 branch_block_stmt_714/ifx_xelse1617_ifx_xend1665_PhiReq/$exit
      -- CP-element group 755: 	 branch_block_stmt_714/ifx_xelse1617_ifx_xend1665_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_755: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_755"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(740) & zeropad3D_CP_2152_elements(748) & zeropad3D_CP_2152_elements(754);
      gj_zeropad3D_cp_element_group_755 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(755), clk => clk, reset => reset); --
    end block;
    -- CP-element group 756:  transition  input  bypass 
    -- CP-element group 756: predecessors 
    -- CP-element group 756: 	1210 
    -- CP-element group 756: successors 
    -- CP-element group 756:  members (3) 
      -- CP-element group 756: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/type_cast_5145_sample_completed_
      -- CP-element group 756: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/type_cast_5145_Sample/$exit
      -- CP-element group 756: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/type_cast_5145_Sample/ra
      -- 
    ra_10769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 756_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5145_inst_ack_0, ack => zeropad3D_CP_2152_elements(756)); -- 
    -- CP-element group 757:  branch  transition  place  input  output  bypass 
    -- CP-element group 757: predecessors 
    -- CP-element group 757: 	1210 
    -- CP-element group 757: successors 
    -- CP-element group 757: 	758 
    -- CP-element group 757: 	759 
    -- CP-element group 757:  members (13) 
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159__exit__
      -- CP-element group 757: 	 branch_block_stmt_714/if_stmt_5160__entry__
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/$exit
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/type_cast_5145_update_completed_
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/type_cast_5145_Update/$exit
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/type_cast_5145_Update/ca
      -- CP-element group 757: 	 branch_block_stmt_714/if_stmt_5160_dead_link/$entry
      -- CP-element group 757: 	 branch_block_stmt_714/if_stmt_5160_eval_test/$entry
      -- CP-element group 757: 	 branch_block_stmt_714/if_stmt_5160_eval_test/$exit
      -- CP-element group 757: 	 branch_block_stmt_714/if_stmt_5160_eval_test/branch_req
      -- CP-element group 757: 	 branch_block_stmt_714/R_cmp1673_5161_place
      -- CP-element group 757: 	 branch_block_stmt_714/if_stmt_5160_if_link/$entry
      -- CP-element group 757: 	 branch_block_stmt_714/if_stmt_5160_else_link/$entry
      -- 
    ca_10774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 757_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5145_inst_ack_1, ack => zeropad3D_CP_2152_elements(757)); -- 
    branch_req_10782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(757), ack => if_stmt_5160_branch_req_0); -- 
    -- CP-element group 758:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 758: predecessors 
    -- CP-element group 758: 	757 
    -- CP-element group 758: successors 
    -- CP-element group 758: 	1219 
    -- CP-element group 758: 	1220 
    -- CP-element group 758: 	1222 
    -- CP-element group 758: 	1223 
    -- CP-element group 758: 	1225 
    -- CP-element group 758: 	1226 
    -- CP-element group 758:  members (40) 
      -- CP-element group 758: 	 branch_block_stmt_714/merge_stmt_5166__exit__
      -- CP-element group 758: 	 branch_block_stmt_714/assign_stmt_5172__entry__
      -- CP-element group 758: 	 branch_block_stmt_714/assign_stmt_5172__exit__
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715
      -- CP-element group 758: 	 branch_block_stmt_714/if_stmt_5160_if_link/$exit
      -- CP-element group 758: 	 branch_block_stmt_714/if_stmt_5160_if_link/if_choice_transition
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xend1665_ifx_xthen1675
      -- CP-element group 758: 	 branch_block_stmt_714/assign_stmt_5172/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/assign_stmt_5172/$exit
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/type_cast_5250/SplitProtocol/Update/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/merge_stmt_5166_PhiReqMerge
      -- CP-element group 758: 	 branch_block_stmt_714/merge_stmt_5166_PhiAck/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/merge_stmt_5166_PhiAck/$exit
      -- CP-element group 758: 	 branch_block_stmt_714/merge_stmt_5166_PhiAck/dummy
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5265/SplitProtocol/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5265/SplitProtocol/Sample/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5265/SplitProtocol/Sample/rr
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/type_cast_5250/SplitProtocol/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xend1665_ifx_xthen1675_PhiReq/$exit
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xend1665_ifx_xthen1675_PhiReq/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/type_cast_5250/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/type_cast_5250/SplitProtocol/Sample/rr
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5265/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5257/SplitProtocol/Update/cr
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5257/SplitProtocol/Update/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5257/SplitProtocol/Sample/rr
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5257/SplitProtocol/Sample/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5257/SplitProtocol/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5257/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5265/SplitProtocol/Update/cr
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5265/SplitProtocol/Update/$entry
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/type_cast_5250/SplitProtocol/Update/cr
      -- CP-element group 758: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/type_cast_5250/SplitProtocol/Sample/$entry
      -- 
    if_choice_transition_10787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 758_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_5160_branch_ack_1, ack => zeropad3D_CP_2152_elements(758)); -- 
    rr_14300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(758), ack => type_cast_5265_inst_req_0); -- 
    rr_14254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(758), ack => type_cast_5250_inst_req_0); -- 
    cr_14282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(758), ack => type_cast_5257_inst_req_1); -- 
    rr_14277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(758), ack => type_cast_5257_inst_req_0); -- 
    cr_14305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(758), ack => type_cast_5265_inst_req_1); -- 
    cr_14259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(758), ack => type_cast_5250_inst_req_1); -- 
    -- CP-element group 759:  fork  transition  place  input  output  bypass 
    -- CP-element group 759: predecessors 
    -- CP-element group 759: 	757 
    -- CP-element group 759: successors 
    -- CP-element group 759: 	760 
    -- CP-element group 759: 	761 
    -- CP-element group 759: 	762 
    -- CP-element group 759: 	763 
    -- CP-element group 759: 	765 
    -- CP-element group 759: 	768 
    -- CP-element group 759: 	770 
    -- CP-element group 759: 	771 
    -- CP-element group 759: 	772 
    -- CP-element group 759: 	774 
    -- CP-element group 759:  members (54) 
      -- CP-element group 759: 	 branch_block_stmt_714/merge_stmt_5174__exit__
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239__entry__
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Sample/word_access_start/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Update/word_access_complete/word_0/cr
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Update/word_access_complete/word_0/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5228_Update/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Update/word_access_complete/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Update/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Sample/word_access_start/word_0/rr
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Sample/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_root_address_calculated
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_word_address_calculated
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_update_start_
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_sample_start_
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5228_update_start_
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5228_Update/cr
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Sample/word_access_start/word_0/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/if_stmt_5160_else_link/$exit
      -- CP-element group 759: 	 branch_block_stmt_714/if_stmt_5160_else_link/else_choice_transition
      -- CP-element group 759: 	 branch_block_stmt_714/ifx_xend1665_ifx_xelse1680
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5184_sample_start_
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5184_update_start_
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5184_Sample/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5184_Sample/rr
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5184_Update/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5184_Update/cr
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_sample_start_
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_update_start_
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_word_address_calculated
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_root_address_calculated
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Sample/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Sample/word_access_start/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Sample/word_access_start/word_0/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Sample/word_access_start/word_0/rr
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Update/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Update/word_access_complete/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Update/word_access_complete/word_0/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Update/word_access_complete/word_0/cr
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5191_update_start_
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5191_Update/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5191_Update/cr
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5205_update_start_
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5205_Update/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5205_Update/cr
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5221_update_start_
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5221_Update/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5221_Update/cr
      -- CP-element group 759: 	 branch_block_stmt_714/ifx_xend1665_ifx_xelse1680_PhiReq/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/ifx_xend1665_ifx_xelse1680_PhiReq/$exit
      -- CP-element group 759: 	 branch_block_stmt_714/merge_stmt_5174_PhiReqMerge
      -- CP-element group 759: 	 branch_block_stmt_714/merge_stmt_5174_PhiAck/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/merge_stmt_5174_PhiAck/$exit
      -- CP-element group 759: 	 branch_block_stmt_714/merge_stmt_5174_PhiAck/dummy
      -- 
    else_choice_transition_10791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 759_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_5160_branch_ack_0, ack => zeropad3D_CP_2152_elements(759)); -- 
    cr_10915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(759), ack => LOAD_row_high_5224_load_0_req_1); -- 
    rr_10904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(759), ack => LOAD_row_high_5224_load_0_req_0); -- 
    cr_10934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(759), ack => type_cast_5228_inst_req_1); -- 
    rr_10807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(759), ack => type_cast_5184_inst_req_0); -- 
    cr_10812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(759), ack => type_cast_5184_inst_req_1); -- 
    rr_10829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(759), ack => LOAD_col_high_5187_load_0_req_0); -- 
    cr_10840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(759), ack => LOAD_col_high_5187_load_0_req_1); -- 
    cr_10859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(759), ack => type_cast_5191_inst_req_1); -- 
    cr_10873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(759), ack => type_cast_5205_inst_req_1); -- 
    cr_10887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(759), ack => type_cast_5221_inst_req_1); -- 
    -- CP-element group 760:  transition  input  bypass 
    -- CP-element group 760: predecessors 
    -- CP-element group 760: 	759 
    -- CP-element group 760: successors 
    -- CP-element group 760:  members (3) 
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5184_sample_completed_
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5184_Sample/$exit
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5184_Sample/ra
      -- 
    ra_10808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 760_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5184_inst_ack_0, ack => zeropad3D_CP_2152_elements(760)); -- 
    -- CP-element group 761:  transition  input  bypass 
    -- CP-element group 761: predecessors 
    -- CP-element group 761: 	759 
    -- CP-element group 761: successors 
    -- CP-element group 761: 	766 
    -- CP-element group 761:  members (3) 
      -- CP-element group 761: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5184_update_completed_
      -- CP-element group 761: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5184_Update/$exit
      -- CP-element group 761: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5184_Update/ca
      -- 
    ca_10813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 761_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5184_inst_ack_1, ack => zeropad3D_CP_2152_elements(761)); -- 
    -- CP-element group 762:  transition  input  bypass 
    -- CP-element group 762: predecessors 
    -- CP-element group 762: 	759 
    -- CP-element group 762: successors 
    -- CP-element group 762:  members (5) 
      -- CP-element group 762: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_sample_completed_
      -- CP-element group 762: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Sample/$exit
      -- CP-element group 762: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Sample/word_access_start/$exit
      -- CP-element group 762: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Sample/word_access_start/word_0/$exit
      -- CP-element group 762: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Sample/word_access_start/word_0/ra
      -- 
    ra_10830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 762_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_5187_load_0_ack_0, ack => zeropad3D_CP_2152_elements(762)); -- 
    -- CP-element group 763:  transition  input  output  bypass 
    -- CP-element group 763: predecessors 
    -- CP-element group 763: 	759 
    -- CP-element group 763: successors 
    -- CP-element group 763: 	764 
    -- CP-element group 763:  members (12) 
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_update_completed_
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Update/$exit
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Update/word_access_complete/$exit
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Update/word_access_complete/word_0/$exit
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Update/word_access_complete/word_0/ca
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Update/LOAD_col_high_5187_Merge/$entry
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Update/LOAD_col_high_5187_Merge/$exit
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Update/LOAD_col_high_5187_Merge/merge_req
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_col_high_5187_Update/LOAD_col_high_5187_Merge/merge_ack
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5191_sample_start_
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5191_Sample/$entry
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5191_Sample/rr
      -- 
    ca_10841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 763_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_5187_load_0_ack_1, ack => zeropad3D_CP_2152_elements(763)); -- 
    rr_10854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(763), ack => type_cast_5191_inst_req_0); -- 
    -- CP-element group 764:  transition  input  bypass 
    -- CP-element group 764: predecessors 
    -- CP-element group 764: 	763 
    -- CP-element group 764: successors 
    -- CP-element group 764:  members (3) 
      -- CP-element group 764: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5191_sample_completed_
      -- CP-element group 764: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5191_Sample/$exit
      -- CP-element group 764: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5191_Sample/ra
      -- 
    ra_10855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 764_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5191_inst_ack_0, ack => zeropad3D_CP_2152_elements(764)); -- 
    -- CP-element group 765:  transition  input  bypass 
    -- CP-element group 765: predecessors 
    -- CP-element group 765: 	759 
    -- CP-element group 765: successors 
    -- CP-element group 765: 	766 
    -- CP-element group 765:  members (3) 
      -- CP-element group 765: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5191_update_completed_
      -- CP-element group 765: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5191_Update/$exit
      -- CP-element group 765: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5191_Update/ca
      -- 
    ca_10860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 765_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5191_inst_ack_1, ack => zeropad3D_CP_2152_elements(765)); -- 
    -- CP-element group 766:  join  transition  output  bypass 
    -- CP-element group 766: predecessors 
    -- CP-element group 766: 	761 
    -- CP-element group 766: 	765 
    -- CP-element group 766: successors 
    -- CP-element group 766: 	767 
    -- CP-element group 766:  members (3) 
      -- CP-element group 766: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5205_sample_start_
      -- CP-element group 766: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5205_Sample/$entry
      -- CP-element group 766: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5205_Sample/rr
      -- 
    rr_10868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(766), ack => type_cast_5205_inst_req_0); -- 
    zeropad3D_cp_element_group_766: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_766"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(761) & zeropad3D_CP_2152_elements(765);
      gj_zeropad3D_cp_element_group_766 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(766), clk => clk, reset => reset); --
    end block;
    -- CP-element group 767:  transition  input  bypass 
    -- CP-element group 767: predecessors 
    -- CP-element group 767: 	766 
    -- CP-element group 767: successors 
    -- CP-element group 767:  members (3) 
      -- CP-element group 767: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5205_sample_completed_
      -- CP-element group 767: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5205_Sample/$exit
      -- CP-element group 767: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5205_Sample/ra
      -- 
    ra_10869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 767_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5205_inst_ack_0, ack => zeropad3D_CP_2152_elements(767)); -- 
    -- CP-element group 768:  transition  input  output  bypass 
    -- CP-element group 768: predecessors 
    -- CP-element group 768: 	759 
    -- CP-element group 768: successors 
    -- CP-element group 768: 	769 
    -- CP-element group 768:  members (6) 
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5205_update_completed_
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5205_Update/$exit
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5205_Update/ca
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5221_sample_start_
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5221_Sample/$entry
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5221_Sample/rr
      -- 
    ca_10874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 768_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5205_inst_ack_1, ack => zeropad3D_CP_2152_elements(768)); -- 
    rr_10882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(768), ack => type_cast_5221_inst_req_0); -- 
    -- CP-element group 769:  transition  input  bypass 
    -- CP-element group 769: predecessors 
    -- CP-element group 769: 	768 
    -- CP-element group 769: successors 
    -- CP-element group 769:  members (3) 
      -- CP-element group 769: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5221_sample_completed_
      -- CP-element group 769: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5221_Sample/$exit
      -- CP-element group 769: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5221_Sample/ra
      -- 
    ra_10883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 769_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5221_inst_ack_0, ack => zeropad3D_CP_2152_elements(769)); -- 
    -- CP-element group 770:  transition  input  bypass 
    -- CP-element group 770: predecessors 
    -- CP-element group 770: 	759 
    -- CP-element group 770: successors 
    -- CP-element group 770: 	775 
    -- CP-element group 770:  members (3) 
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5221_Update/ca
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5221_update_completed_
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5221_Update/$exit
      -- 
    ca_10888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 770_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5221_inst_ack_1, ack => zeropad3D_CP_2152_elements(770)); -- 
    -- CP-element group 771:  transition  input  bypass 
    -- CP-element group 771: predecessors 
    -- CP-element group 771: 	759 
    -- CP-element group 771: successors 
    -- CP-element group 771:  members (5) 
      -- CP-element group 771: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Sample/word_access_start/$exit
      -- CP-element group 771: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Sample/$exit
      -- CP-element group 771: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Sample/word_access_start/word_0/ra
      -- CP-element group 771: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Sample/word_access_start/word_0/$exit
      -- CP-element group 771: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_sample_completed_
      -- 
    ra_10905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 771_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_5224_load_0_ack_0, ack => zeropad3D_CP_2152_elements(771)); -- 
    -- CP-element group 772:  transition  input  output  bypass 
    -- CP-element group 772: predecessors 
    -- CP-element group 772: 	759 
    -- CP-element group 772: successors 
    -- CP-element group 772: 	773 
    -- CP-element group 772:  members (12) 
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Update/LOAD_row_high_5224_Merge/merge_req
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Update/LOAD_row_high_5224_Merge/$exit
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Update/LOAD_row_high_5224_Merge/$entry
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Update/word_access_complete/word_0/ca
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Update/word_access_complete/word_0/$exit
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Update/word_access_complete/$exit
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Update/$exit
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5228_Sample/rr
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_update_completed_
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5228_Sample/$entry
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5228_sample_start_
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/LOAD_row_high_5224_Update/LOAD_row_high_5224_Merge/merge_ack
      -- 
    ca_10916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 772_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_5224_load_0_ack_1, ack => zeropad3D_CP_2152_elements(772)); -- 
    rr_10929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(772), ack => type_cast_5228_inst_req_0); -- 
    -- CP-element group 773:  transition  input  bypass 
    -- CP-element group 773: predecessors 
    -- CP-element group 773: 	772 
    -- CP-element group 773: successors 
    -- CP-element group 773:  members (3) 
      -- CP-element group 773: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5228_Sample/ra
      -- CP-element group 773: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5228_Sample/$exit
      -- CP-element group 773: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5228_sample_completed_
      -- 
    ra_10930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 773_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5228_inst_ack_0, ack => zeropad3D_CP_2152_elements(773)); -- 
    -- CP-element group 774:  transition  input  bypass 
    -- CP-element group 774: predecessors 
    -- CP-element group 774: 	759 
    -- CP-element group 774: successors 
    -- CP-element group 774: 	775 
    -- CP-element group 774:  members (3) 
      -- CP-element group 774: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5228_Update/$exit
      -- CP-element group 774: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5228_Update/ca
      -- CP-element group 774: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/type_cast_5228_update_completed_
      -- 
    ca_10935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 774_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5228_inst_ack_1, ack => zeropad3D_CP_2152_elements(774)); -- 
    -- CP-element group 775:  branch  join  transition  place  output  bypass 
    -- CP-element group 775: predecessors 
    -- CP-element group 775: 	770 
    -- CP-element group 775: 	774 
    -- CP-element group 775: successors 
    -- CP-element group 775: 	776 
    -- CP-element group 775: 	777 
    -- CP-element group 775:  members (10) 
      -- CP-element group 775: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239__exit__
      -- CP-element group 775: 	 branch_block_stmt_714/if_stmt_5240__entry__
      -- CP-element group 775: 	 branch_block_stmt_714/if_stmt_5240_if_link/$entry
      -- CP-element group 775: 	 branch_block_stmt_714/if_stmt_5240_eval_test/branch_req
      -- CP-element group 775: 	 branch_block_stmt_714/if_stmt_5240_eval_test/$exit
      -- CP-element group 775: 	 branch_block_stmt_714/if_stmt_5240_eval_test/$entry
      -- CP-element group 775: 	 branch_block_stmt_714/R_cmp1706_5241_place
      -- CP-element group 775: 	 branch_block_stmt_714/if_stmt_5240_dead_link/$entry
      -- CP-element group 775: 	 branch_block_stmt_714/if_stmt_5240_else_link/$entry
      -- CP-element group 775: 	 branch_block_stmt_714/assign_stmt_5180_to_assign_stmt_5239/$exit
      -- 
    branch_req_10943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(775), ack => if_stmt_5240_branch_req_0); -- 
    zeropad3D_cp_element_group_775: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_775"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(770) & zeropad3D_CP_2152_elements(774);
      gj_zeropad3D_cp_element_group_775 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(775), clk => clk, reset => reset); --
    end block;
    -- CP-element group 776:  fork  transition  place  input  output  bypass 
    -- CP-element group 776: predecessors 
    -- CP-element group 776: 	775 
    -- CP-element group 776: successors 
    -- CP-element group 776: 	778 
    -- CP-element group 776: 	779 
    -- CP-element group 776:  members (18) 
      -- CP-element group 776: 	 branch_block_stmt_714/merge_stmt_5268__exit__
      -- CP-element group 776: 	 branch_block_stmt_714/call_stmt_5270__entry__
      -- CP-element group 776: 	 branch_block_stmt_714/if_stmt_5240_if_link/$exit
      -- CP-element group 776: 	 branch_block_stmt_714/ifx_xelse1680_whilex_xend1716
      -- CP-element group 776: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Update/ccr
      -- CP-element group 776: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Update/$entry
      -- CP-element group 776: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Sample/crr
      -- CP-element group 776: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Sample/$entry
      -- CP-element group 776: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_update_start_
      -- CP-element group 776: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_sample_start_
      -- CP-element group 776: 	 branch_block_stmt_714/call_stmt_5270/$entry
      -- CP-element group 776: 	 branch_block_stmt_714/if_stmt_5240_if_link/if_choice_transition
      -- CP-element group 776: 	 branch_block_stmt_714/ifx_xelse1680_whilex_xend1716_PhiReq/$entry
      -- CP-element group 776: 	 branch_block_stmt_714/ifx_xelse1680_whilex_xend1716_PhiReq/$exit
      -- CP-element group 776: 	 branch_block_stmt_714/merge_stmt_5268_PhiReqMerge
      -- CP-element group 776: 	 branch_block_stmt_714/merge_stmt_5268_PhiAck/$entry
      -- CP-element group 776: 	 branch_block_stmt_714/merge_stmt_5268_PhiAck/$exit
      -- CP-element group 776: 	 branch_block_stmt_714/merge_stmt_5268_PhiAck/dummy
      -- 
    if_choice_transition_10948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 776_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_5240_branch_ack_1, ack => zeropad3D_CP_2152_elements(776)); -- 
    ccr_10970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_10970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(776), ack => call_stmt_5270_call_req_1); -- 
    crr_10965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_10965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(776), ack => call_stmt_5270_call_req_0); -- 
    -- CP-element group 777:  fork  transition  place  input  output  bypass 
    -- CP-element group 777: predecessors 
    -- CP-element group 777: 	775 
    -- CP-element group 777: successors 
    -- CP-element group 777: 	1211 
    -- CP-element group 777: 	1212 
    -- CP-element group 777: 	1213 
    -- CP-element group 777: 	1215 
    -- CP-element group 777: 	1216 
    -- CP-element group 777:  members (22) 
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715
      -- CP-element group 777: 	 branch_block_stmt_714/if_stmt_5240_else_link/else_choice_transition
      -- CP-element group 777: 	 branch_block_stmt_714/if_stmt_5240_else_link/$exit
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5263/SplitProtocol/Sample/rr
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5263/SplitProtocol/Update/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5263/SplitProtocol/Update/cr
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5263/SplitProtocol/Sample/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5263/SplitProtocol/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5263/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5259/SplitProtocol/Update/cr
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5247/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5259/SplitProtocol/Update/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5259/SplitProtocol/Sample/rr
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5259/SplitProtocol/Sample/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5259/SplitProtocol/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5259/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/$entry
      -- 
    else_choice_transition_10952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 777_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_5240_branch_ack_0, ack => zeropad3D_CP_2152_elements(777)); -- 
    rr_14228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(777), ack => type_cast_5263_inst_req_0); -- 
    cr_14233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(777), ack => type_cast_5263_inst_req_1); -- 
    cr_14210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(777), ack => type_cast_5259_inst_req_1); -- 
    rr_14205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(777), ack => type_cast_5259_inst_req_0); -- 
    -- CP-element group 778:  transition  input  bypass 
    -- CP-element group 778: predecessors 
    -- CP-element group 778: 	776 
    -- CP-element group 778: successors 
    -- CP-element group 778:  members (3) 
      -- CP-element group 778: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Sample/cra
      -- CP-element group 778: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Sample/$exit
      -- CP-element group 778: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_sample_completed_
      -- 
    cra_10966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 778_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_5270_call_ack_0, ack => zeropad3D_CP_2152_elements(778)); -- 
    -- CP-element group 779:  transition  place  input  bypass 
    -- CP-element group 779: predecessors 
    -- CP-element group 779: 	776 
    -- CP-element group 779: successors 
    -- CP-element group 779:  members (16) 
      -- CP-element group 779: 	 branch_block_stmt_714/branch_block_stmt_714__exit__
      -- CP-element group 779: 	 branch_block_stmt_714/$exit
      -- CP-element group 779: 	 $exit
      -- CP-element group 779: 	 branch_block_stmt_714/call_stmt_5270__exit__
      -- CP-element group 779: 	 branch_block_stmt_714/return__
      -- CP-element group 779: 	 branch_block_stmt_714/merge_stmt_5272__exit__
      -- CP-element group 779: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Update/cca
      -- CP-element group 779: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Update/$exit
      -- CP-element group 779: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_update_completed_
      -- CP-element group 779: 	 branch_block_stmt_714/call_stmt_5270/$exit
      -- CP-element group 779: 	 branch_block_stmt_714/return___PhiReq/$entry
      -- CP-element group 779: 	 branch_block_stmt_714/return___PhiReq/$exit
      -- CP-element group 779: 	 branch_block_stmt_714/merge_stmt_5272_PhiReqMerge
      -- CP-element group 779: 	 branch_block_stmt_714/merge_stmt_5272_PhiAck/$entry
      -- CP-element group 779: 	 branch_block_stmt_714/merge_stmt_5272_PhiAck/$exit
      -- CP-element group 779: 	 branch_block_stmt_714/merge_stmt_5272_PhiAck/dummy
      -- 
    cca_10971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 779_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_5270_call_ack_1, ack => zeropad3D_CP_2152_elements(779)); -- 
    -- CP-element group 780:  transition  output  delay-element  bypass 
    -- CP-element group 780: predecessors 
    -- CP-element group 780: 	58 
    -- CP-element group 780: successors 
    -- CP-element group 780: 	783 
    -- CP-element group 780:  members (4) 
      -- CP-element group 780: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_req
      -- CP-element group 780: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_903_konst_delay_trans
      -- CP-element group 780: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/$exit
      -- CP-element group 780: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_899/$exit
      -- 
    phi_stmt_899_req_10982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_899_req_10982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(780), ack => phi_stmt_899_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(780) is a control-delay.
    cp_element_780_delay: control_delay_element  generic map(name => " 780_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(58), ack => zeropad3D_CP_2152_elements(780), clk => clk, reset =>reset);
    -- CP-element group 781:  transition  output  delay-element  bypass 
    -- CP-element group 781: predecessors 
    -- CP-element group 781: 	58 
    -- CP-element group 781: successors 
    -- CP-element group 781: 	783 
    -- CP-element group 781:  members (4) 
      -- CP-element group 781: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_req
      -- CP-element group 781: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_910_konst_delay_trans
      -- CP-element group 781: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/$exit
      -- CP-element group 781: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_906/$exit
      -- 
    phi_stmt_906_req_10990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_906_req_10990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(781), ack => phi_stmt_906_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(781) is a control-delay.
    cp_element_781_delay: control_delay_element  generic map(name => " 781_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(58), ack => zeropad3D_CP_2152_elements(781), clk => clk, reset =>reset);
    -- CP-element group 782:  transition  output  delay-element  bypass 
    -- CP-element group 782: predecessors 
    -- CP-element group 782: 	58 
    -- CP-element group 782: successors 
    -- CP-element group 782: 	783 
    -- CP-element group 782:  members (4) 
      -- CP-element group 782: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_req
      -- CP-element group 782: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_917_konst_delay_trans
      -- CP-element group 782: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/$exit
      -- CP-element group 782: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_913/$exit
      -- 
    phi_stmt_913_req_10998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_913_req_10998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(782), ack => phi_stmt_913_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(782) is a control-delay.
    cp_element_782_delay: control_delay_element  generic map(name => " 782_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(58), ack => zeropad3D_CP_2152_elements(782), clk => clk, reset =>reset);
    -- CP-element group 783:  join  transition  bypass 
    -- CP-element group 783: predecessors 
    -- CP-element group 783: 	780 
    -- CP-element group 783: 	781 
    -- CP-element group 783: 	782 
    -- CP-element group 783: successors 
    -- CP-element group 783: 	794 
    -- CP-element group 783:  members (1) 
      -- CP-element group 783: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_783: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_783"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(780) & zeropad3D_CP_2152_elements(781) & zeropad3D_CP_2152_elements(782);
      gj_zeropad3D_cp_element_group_783 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(783), clk => clk, reset => reset); --
    end block;
    -- CP-element group 784:  transition  input  bypass 
    -- CP-element group 784: predecessors 
    -- CP-element group 784: 	1 
    -- CP-element group 784: successors 
    -- CP-element group 784: 	786 
    -- CP-element group 784:  members (2) 
      -- CP-element group 784: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Sample/ra
      -- CP-element group 784: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Sample/$exit
      -- 
    ra_11018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 784_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_0, ack => zeropad3D_CP_2152_elements(784)); -- 
    -- CP-element group 785:  transition  input  bypass 
    -- CP-element group 785: predecessors 
    -- CP-element group 785: 	1 
    -- CP-element group 785: successors 
    -- CP-element group 785: 	786 
    -- CP-element group 785:  members (2) 
      -- CP-element group 785: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Update/ca
      -- CP-element group 785: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Update/$exit
      -- 
    ca_11023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 785_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_1, ack => zeropad3D_CP_2152_elements(785)); -- 
    -- CP-element group 786:  join  transition  output  bypass 
    -- CP-element group 786: predecessors 
    -- CP-element group 786: 	784 
    -- CP-element group 786: 	785 
    -- CP-element group 786: successors 
    -- CP-element group 786: 	793 
    -- CP-element group 786:  members (5) 
      -- CP-element group 786: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_req
      -- CP-element group 786: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/$exit
      -- CP-element group 786: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/$exit
      -- CP-element group 786: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/$exit
      -- CP-element group 786: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/$exit
      -- 
    phi_stmt_899_req_11024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_899_req_11024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(786), ack => phi_stmt_899_req_1); -- 
    zeropad3D_cp_element_group_786: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_786"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(784) & zeropad3D_CP_2152_elements(785);
      gj_zeropad3D_cp_element_group_786 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(786), clk => clk, reset => reset); --
    end block;
    -- CP-element group 787:  transition  input  bypass 
    -- CP-element group 787: predecessors 
    -- CP-element group 787: 	1 
    -- CP-element group 787: successors 
    -- CP-element group 787: 	789 
    -- CP-element group 787:  members (2) 
      -- CP-element group 787: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Sample/ra
      -- CP-element group 787: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Sample/$exit
      -- 
    ra_11041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 787_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_912_inst_ack_0, ack => zeropad3D_CP_2152_elements(787)); -- 
    -- CP-element group 788:  transition  input  bypass 
    -- CP-element group 788: predecessors 
    -- CP-element group 788: 	1 
    -- CP-element group 788: successors 
    -- CP-element group 788: 	789 
    -- CP-element group 788:  members (2) 
      -- CP-element group 788: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Update/ca
      -- CP-element group 788: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Update/$exit
      -- 
    ca_11046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 788_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_912_inst_ack_1, ack => zeropad3D_CP_2152_elements(788)); -- 
    -- CP-element group 789:  join  transition  output  bypass 
    -- CP-element group 789: predecessors 
    -- CP-element group 789: 	787 
    -- CP-element group 789: 	788 
    -- CP-element group 789: successors 
    -- CP-element group 789: 	793 
    -- CP-element group 789:  members (5) 
      -- CP-element group 789: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/$exit
      -- CP-element group 789: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_req
      -- CP-element group 789: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/$exit
      -- CP-element group 789: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/$exit
      -- CP-element group 789: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/$exit
      -- 
    phi_stmt_906_req_11047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_906_req_11047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(789), ack => phi_stmt_906_req_1); -- 
    zeropad3D_cp_element_group_789: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_789"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(787) & zeropad3D_CP_2152_elements(788);
      gj_zeropad3D_cp_element_group_789 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(789), clk => clk, reset => reset); --
    end block;
    -- CP-element group 790:  transition  input  bypass 
    -- CP-element group 790: predecessors 
    -- CP-element group 790: 	1 
    -- CP-element group 790: successors 
    -- CP-element group 790: 	792 
    -- CP-element group 790:  members (2) 
      -- CP-element group 790: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Sample/ra
      -- CP-element group 790: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Sample/$exit
      -- 
    ra_11064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 790_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_919_inst_ack_0, ack => zeropad3D_CP_2152_elements(790)); -- 
    -- CP-element group 791:  transition  input  bypass 
    -- CP-element group 791: predecessors 
    -- CP-element group 791: 	1 
    -- CP-element group 791: successors 
    -- CP-element group 791: 	792 
    -- CP-element group 791:  members (2) 
      -- CP-element group 791: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Update/ca
      -- CP-element group 791: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Update/$exit
      -- 
    ca_11069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 791_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_919_inst_ack_1, ack => zeropad3D_CP_2152_elements(791)); -- 
    -- CP-element group 792:  join  transition  output  bypass 
    -- CP-element group 792: predecessors 
    -- CP-element group 792: 	790 
    -- CP-element group 792: 	791 
    -- CP-element group 792: successors 
    -- CP-element group 792: 	793 
    -- CP-element group 792:  members (5) 
      -- CP-element group 792: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/$exit
      -- CP-element group 792: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/$exit
      -- CP-element group 792: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_req
      -- CP-element group 792: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/$exit
      -- CP-element group 792: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/$exit
      -- 
    phi_stmt_913_req_11070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_913_req_11070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(792), ack => phi_stmt_913_req_1); -- 
    zeropad3D_cp_element_group_792: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_792"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(790) & zeropad3D_CP_2152_elements(791);
      gj_zeropad3D_cp_element_group_792 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(792), clk => clk, reset => reset); --
    end block;
    -- CP-element group 793:  join  transition  bypass 
    -- CP-element group 793: predecessors 
    -- CP-element group 793: 	786 
    -- CP-element group 793: 	789 
    -- CP-element group 793: 	792 
    -- CP-element group 793: successors 
    -- CP-element group 793: 	794 
    -- CP-element group 793:  members (1) 
      -- CP-element group 793: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_793: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_793"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(786) & zeropad3D_CP_2152_elements(789) & zeropad3D_CP_2152_elements(792);
      gj_zeropad3D_cp_element_group_793 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(793), clk => clk, reset => reset); --
    end block;
    -- CP-element group 794:  merge  fork  transition  place  bypass 
    -- CP-element group 794: predecessors 
    -- CP-element group 794: 	783 
    -- CP-element group 794: 	793 
    -- CP-element group 794: successors 
    -- CP-element group 794: 	795 
    -- CP-element group 794: 	796 
    -- CP-element group 794: 	797 
    -- CP-element group 794:  members (2) 
      -- CP-element group 794: 	 branch_block_stmt_714/merge_stmt_898_PhiReqMerge
      -- CP-element group 794: 	 branch_block_stmt_714/merge_stmt_898_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(794) <= OrReduce(zeropad3D_CP_2152_elements(783) & zeropad3D_CP_2152_elements(793));
    -- CP-element group 795:  transition  input  bypass 
    -- CP-element group 795: predecessors 
    -- CP-element group 795: 	794 
    -- CP-element group 795: successors 
    -- CP-element group 795: 	798 
    -- CP-element group 795:  members (1) 
      -- CP-element group 795: 	 branch_block_stmt_714/merge_stmt_898_PhiAck/phi_stmt_899_ack
      -- 
    phi_stmt_899_ack_11075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 795_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_899_ack_0, ack => zeropad3D_CP_2152_elements(795)); -- 
    -- CP-element group 796:  transition  input  bypass 
    -- CP-element group 796: predecessors 
    -- CP-element group 796: 	794 
    -- CP-element group 796: successors 
    -- CP-element group 796: 	798 
    -- CP-element group 796:  members (1) 
      -- CP-element group 796: 	 branch_block_stmt_714/merge_stmt_898_PhiAck/phi_stmt_906_ack
      -- 
    phi_stmt_906_ack_11076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 796_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_906_ack_0, ack => zeropad3D_CP_2152_elements(796)); -- 
    -- CP-element group 797:  transition  input  bypass 
    -- CP-element group 797: predecessors 
    -- CP-element group 797: 	794 
    -- CP-element group 797: successors 
    -- CP-element group 797: 	798 
    -- CP-element group 797:  members (1) 
      -- CP-element group 797: 	 branch_block_stmt_714/merge_stmt_898_PhiAck/phi_stmt_913_ack
      -- 
    phi_stmt_913_ack_11077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 797_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_913_ack_0, ack => zeropad3D_CP_2152_elements(797)); -- 
    -- CP-element group 798:  join  fork  transition  place  output  bypass 
    -- CP-element group 798: predecessors 
    -- CP-element group 798: 	795 
    -- CP-element group 798: 	796 
    -- CP-element group 798: 	797 
    -- CP-element group 798: successors 
    -- CP-element group 798: 	59 
    -- CP-element group 798: 	60 
    -- CP-element group 798:  members (10) 
      -- CP-element group 798: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932__entry__
      -- CP-element group 798: 	 branch_block_stmt_714/merge_stmt_898__exit__
      -- CP-element group 798: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_sample_start_
      -- CP-element group 798: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_update_start_
      -- CP-element group 798: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Sample/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Sample/rr
      -- CP-element group 798: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Update/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Update/cr
      -- CP-element group 798: 	 branch_block_stmt_714/merge_stmt_898_PhiAck/$exit
      -- 
    rr_3166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(798), ack => type_cast_924_inst_req_0); -- 
    cr_3171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(798), ack => type_cast_924_inst_req_1); -- 
    zeropad3D_cp_element_group_798: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_798"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(795) & zeropad3D_CP_2152_elements(796) & zeropad3D_CP_2152_elements(797);
      gj_zeropad3D_cp_element_group_798 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(798), clk => clk, reset => reset); --
    end block;
    -- CP-element group 799:  merge  fork  transition  place  output  bypass 
    -- CP-element group 799: predecessors 
    -- CP-element group 799: 	61 
    -- CP-element group 799: 	68 
    -- CP-element group 799: 	71 
    -- CP-element group 799: 	78 
    -- CP-element group 799: successors 
    -- CP-element group 799: 	79 
    -- CP-element group 799: 	80 
    -- CP-element group 799: 	81 
    -- CP-element group 799: 	82 
    -- CP-element group 799: 	85 
    -- CP-element group 799: 	87 
    -- CP-element group 799: 	89 
    -- CP-element group 799: 	91 
    -- CP-element group 799:  members (33) 
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079__entry__
      -- CP-element group 799: 	 branch_block_stmt_714/merge_stmt_1022__exit__
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_sample_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Update/cr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_update_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Update/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_update_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_complete/req
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Update/cr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Update/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Sample/rr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_complete/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Sample/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_update_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_update_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/word_access_complete/word_0/cr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Update/req
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Update/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_sample_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/word_access_complete/word_0/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_update_start
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Update/cr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Update/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/word_access_complete/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Sample/rr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Sample/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_update_start_
      -- CP-element group 799: 	 branch_block_stmt_714/merge_stmt_1022_PhiAck/dummy
      -- CP-element group 799: 	 branch_block_stmt_714/merge_stmt_1022_PhiAck/$exit
      -- CP-element group 799: 	 branch_block_stmt_714/merge_stmt_1022_PhiAck/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/merge_stmt_1022_PhiReqMerge
      -- 
    cr_3381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => type_cast_1026_inst_req_1); -- 
    req_3455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => addr_of_1073_final_reg_req_1); -- 
    cr_3409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => type_cast_1066_inst_req_1); -- 
    rr_3376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => type_cast_1026_inst_req_0); -- 
    cr_3505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => ptr_deref_1076_store_0_req_1); -- 
    req_3440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => array_obj_ref_1072_index_offset_req_1); -- 
    cr_3395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => type_cast_1031_inst_req_1); -- 
    rr_3390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => type_cast_1031_inst_req_0); -- 
    zeropad3D_CP_2152_elements(799) <= OrReduce(zeropad3D_CP_2152_elements(61) & zeropad3D_CP_2152_elements(68) & zeropad3D_CP_2152_elements(71) & zeropad3D_CP_2152_elements(78));
    -- CP-element group 800:  merge  fork  transition  place  output  bypass 
    -- CP-element group 800: predecessors 
    -- CP-element group 800: 	92 
    -- CP-element group 800: 	112 
    -- CP-element group 800: successors 
    -- CP-element group 800: 	113 
    -- CP-element group 800: 	114 
    -- CP-element group 800:  members (13) 
      -- CP-element group 800: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206__entry__
      -- CP-element group 800: 	 branch_block_stmt_714/merge_stmt_1188__exit__
      -- CP-element group 800: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/$entry
      -- CP-element group 800: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_sample_start_
      -- CP-element group 800: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_update_start_
      -- CP-element group 800: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Sample/$entry
      -- CP-element group 800: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Sample/rr
      -- CP-element group 800: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Update/$entry
      -- CP-element group 800: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Update/cr
      -- CP-element group 800: 	 branch_block_stmt_714/merge_stmt_1188_PhiAck/dummy
      -- CP-element group 800: 	 branch_block_stmt_714/merge_stmt_1188_PhiAck/$exit
      -- CP-element group 800: 	 branch_block_stmt_714/merge_stmt_1188_PhiAck/$entry
      -- CP-element group 800: 	 branch_block_stmt_714/merge_stmt_1188_PhiReqMerge
      -- 
    rr_3754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(800), ack => type_cast_1192_inst_req_0); -- 
    cr_3759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(800), ack => type_cast_1192_inst_req_1); -- 
    zeropad3D_CP_2152_elements(800) <= OrReduce(zeropad3D_CP_2152_elements(92) & zeropad3D_CP_2152_elements(112));
    -- CP-element group 801:  transition  input  bypass 
    -- CP-element group 801: predecessors 
    -- CP-element group 801: 	134 
    -- CP-element group 801: successors 
    -- CP-element group 801: 	803 
    -- CP-element group 801:  members (2) 
      -- CP-element group 801: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Sample/$exit
      -- CP-element group 801: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Sample/ra
      -- 
    ra_11197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 801_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1318_inst_ack_0, ack => zeropad3D_CP_2152_elements(801)); -- 
    -- CP-element group 802:  transition  input  bypass 
    -- CP-element group 802: predecessors 
    -- CP-element group 802: 	134 
    -- CP-element group 802: successors 
    -- CP-element group 802: 	803 
    -- CP-element group 802:  members (2) 
      -- CP-element group 802: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Update/$exit
      -- CP-element group 802: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Update/ca
      -- 
    ca_11202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 802_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1318_inst_ack_1, ack => zeropad3D_CP_2152_elements(802)); -- 
    -- CP-element group 803:  join  transition  output  bypass 
    -- CP-element group 803: predecessors 
    -- CP-element group 803: 	801 
    -- CP-element group 803: 	802 
    -- CP-element group 803: successors 
    -- CP-element group 803: 	808 
    -- CP-element group 803:  members (5) 
      -- CP-element group 803: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/$exit
      -- CP-element group 803: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/$exit
      -- CP-element group 803: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/$exit
      -- CP-element group 803: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_req
      -- CP-element group 803: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/$exit
      -- 
    phi_stmt_1313_req_11203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1313_req_11203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(803), ack => phi_stmt_1313_req_1); -- 
    zeropad3D_cp_element_group_803: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_803"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(801) & zeropad3D_CP_2152_elements(802);
      gj_zeropad3D_cp_element_group_803 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(803), clk => clk, reset => reset); --
    end block;
    -- CP-element group 804:  transition  output  delay-element  bypass 
    -- CP-element group 804: predecessors 
    -- CP-element group 804: 	134 
    -- CP-element group 804: successors 
    -- CP-element group 804: 	808 
    -- CP-element group 804:  members (4) 
      -- CP-element group 804: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_req
      -- CP-element group 804: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1323_konst_delay_trans
      -- CP-element group 804: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/$exit
      -- CP-element group 804: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1319/$exit
      -- 
    phi_stmt_1319_req_11211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1319_req_11211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(804), ack => phi_stmt_1319_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(804) is a control-delay.
    cp_element_804_delay: control_delay_element  generic map(name => " 804_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(134), ack => zeropad3D_CP_2152_elements(804), clk => clk, reset =>reset);
    -- CP-element group 805:  transition  input  bypass 
    -- CP-element group 805: predecessors 
    -- CP-element group 805: 	134 
    -- CP-element group 805: successors 
    -- CP-element group 805: 	807 
    -- CP-element group 805:  members (2) 
      -- CP-element group 805: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Sample/ra
      -- CP-element group 805: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Sample/$exit
      -- 
    ra_11228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 805_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1310_inst_ack_0, ack => zeropad3D_CP_2152_elements(805)); -- 
    -- CP-element group 806:  transition  input  bypass 
    -- CP-element group 806: predecessors 
    -- CP-element group 806: 	134 
    -- CP-element group 806: successors 
    -- CP-element group 806: 	807 
    -- CP-element group 806:  members (2) 
      -- CP-element group 806: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Update/ca
      -- CP-element group 806: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Update/$exit
      -- 
    ca_11233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 806_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1310_inst_ack_1, ack => zeropad3D_CP_2152_elements(806)); -- 
    -- CP-element group 807:  join  transition  output  bypass 
    -- CP-element group 807: predecessors 
    -- CP-element group 807: 	805 
    -- CP-element group 807: 	806 
    -- CP-element group 807: successors 
    -- CP-element group 807: 	808 
    -- CP-element group 807:  members (5) 
      -- CP-element group 807: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_req
      -- CP-element group 807: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/$exit
      -- CP-element group 807: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/$exit
      -- CP-element group 807: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/$exit
      -- CP-element group 807: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/$exit
      -- 
    phi_stmt_1307_req_11234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1307_req_11234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(807), ack => phi_stmt_1307_req_0); -- 
    zeropad3D_cp_element_group_807: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_807"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(805) & zeropad3D_CP_2152_elements(806);
      gj_zeropad3D_cp_element_group_807 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(807), clk => clk, reset => reset); --
    end block;
    -- CP-element group 808:  join  transition  bypass 
    -- CP-element group 808: predecessors 
    -- CP-element group 808: 	803 
    -- CP-element group 808: 	804 
    -- CP-element group 808: 	807 
    -- CP-element group 808: successors 
    -- CP-element group 808: 	819 
    -- CP-element group 808:  members (1) 
      -- CP-element group 808: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_808: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_808"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(803) & zeropad3D_CP_2152_elements(804) & zeropad3D_CP_2152_elements(807);
      gj_zeropad3D_cp_element_group_808 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(808), clk => clk, reset => reset); --
    end block;
    -- CP-element group 809:  transition  input  bypass 
    -- CP-element group 809: predecessors 
    -- CP-element group 809: 	115 
    -- CP-element group 809: successors 
    -- CP-element group 809: 	811 
    -- CP-element group 809:  members (2) 
      -- CP-element group 809: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Sample/$exit
      -- CP-element group 809: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Sample/ra
      -- 
    ra_11254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 809_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1316_inst_ack_0, ack => zeropad3D_CP_2152_elements(809)); -- 
    -- CP-element group 810:  transition  input  bypass 
    -- CP-element group 810: predecessors 
    -- CP-element group 810: 	115 
    -- CP-element group 810: successors 
    -- CP-element group 810: 	811 
    -- CP-element group 810:  members (2) 
      -- CP-element group 810: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Update/ca
      -- CP-element group 810: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Update/$exit
      -- 
    ca_11259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 810_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1316_inst_ack_1, ack => zeropad3D_CP_2152_elements(810)); -- 
    -- CP-element group 811:  join  transition  output  bypass 
    -- CP-element group 811: predecessors 
    -- CP-element group 811: 	809 
    -- CP-element group 811: 	810 
    -- CP-element group 811: successors 
    -- CP-element group 811: 	818 
    -- CP-element group 811:  members (5) 
      -- CP-element group 811: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/$exit
      -- CP-element group 811: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/$exit
      -- CP-element group 811: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/$exit
      -- CP-element group 811: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/$exit
      -- CP-element group 811: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_req
      -- 
    phi_stmt_1313_req_11260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1313_req_11260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(811), ack => phi_stmt_1313_req_0); -- 
    zeropad3D_cp_element_group_811: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_811"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(809) & zeropad3D_CP_2152_elements(810);
      gj_zeropad3D_cp_element_group_811 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(811), clk => clk, reset => reset); --
    end block;
    -- CP-element group 812:  transition  input  bypass 
    -- CP-element group 812: predecessors 
    -- CP-element group 812: 	115 
    -- CP-element group 812: successors 
    -- CP-element group 812: 	814 
    -- CP-element group 812:  members (2) 
      -- CP-element group 812: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Sample/$exit
      -- CP-element group 812: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Sample/ra
      -- 
    ra_11277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 812_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1325_inst_ack_0, ack => zeropad3D_CP_2152_elements(812)); -- 
    -- CP-element group 813:  transition  input  bypass 
    -- CP-element group 813: predecessors 
    -- CP-element group 813: 	115 
    -- CP-element group 813: successors 
    -- CP-element group 813: 	814 
    -- CP-element group 813:  members (2) 
      -- CP-element group 813: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Update/ca
      -- CP-element group 813: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Update/$exit
      -- 
    ca_11282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 813_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1325_inst_ack_1, ack => zeropad3D_CP_2152_elements(813)); -- 
    -- CP-element group 814:  join  transition  output  bypass 
    -- CP-element group 814: predecessors 
    -- CP-element group 814: 	812 
    -- CP-element group 814: 	813 
    -- CP-element group 814: successors 
    -- CP-element group 814: 	818 
    -- CP-element group 814:  members (5) 
      -- CP-element group 814: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/$exit
      -- CP-element group 814: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/$exit
      -- CP-element group 814: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/$exit
      -- CP-element group 814: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/$exit
      -- CP-element group 814: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_req
      -- 
    phi_stmt_1319_req_11283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1319_req_11283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(814), ack => phi_stmt_1319_req_1); -- 
    zeropad3D_cp_element_group_814: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_814"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(812) & zeropad3D_CP_2152_elements(813);
      gj_zeropad3D_cp_element_group_814 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(814), clk => clk, reset => reset); --
    end block;
    -- CP-element group 815:  transition  input  bypass 
    -- CP-element group 815: predecessors 
    -- CP-element group 815: 	115 
    -- CP-element group 815: successors 
    -- CP-element group 815: 	817 
    -- CP-element group 815:  members (2) 
      -- CP-element group 815: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Sample/ra
      -- CP-element group 815: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Sample/$exit
      -- 
    ra_11300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 815_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1312_inst_ack_0, ack => zeropad3D_CP_2152_elements(815)); -- 
    -- CP-element group 816:  transition  input  bypass 
    -- CP-element group 816: predecessors 
    -- CP-element group 816: 	115 
    -- CP-element group 816: successors 
    -- CP-element group 816: 	817 
    -- CP-element group 816:  members (2) 
      -- CP-element group 816: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Update/ca
      -- CP-element group 816: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Update/$exit
      -- 
    ca_11305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 816_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1312_inst_ack_1, ack => zeropad3D_CP_2152_elements(816)); -- 
    -- CP-element group 817:  join  transition  output  bypass 
    -- CP-element group 817: predecessors 
    -- CP-element group 817: 	815 
    -- CP-element group 817: 	816 
    -- CP-element group 817: successors 
    -- CP-element group 817: 	818 
    -- CP-element group 817:  members (5) 
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/$exit
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/$exit
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/$exit
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/$exit
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_req
      -- 
    phi_stmt_1307_req_11306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1307_req_11306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(817), ack => phi_stmt_1307_req_1); -- 
    zeropad3D_cp_element_group_817: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_817"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(815) & zeropad3D_CP_2152_elements(816);
      gj_zeropad3D_cp_element_group_817 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(817), clk => clk, reset => reset); --
    end block;
    -- CP-element group 818:  join  transition  bypass 
    -- CP-element group 818: predecessors 
    -- CP-element group 818: 	811 
    -- CP-element group 818: 	814 
    -- CP-element group 818: 	817 
    -- CP-element group 818: successors 
    -- CP-element group 818: 	819 
    -- CP-element group 818:  members (1) 
      -- CP-element group 818: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_818: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_818"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(811) & zeropad3D_CP_2152_elements(814) & zeropad3D_CP_2152_elements(817);
      gj_zeropad3D_cp_element_group_818 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(818), clk => clk, reset => reset); --
    end block;
    -- CP-element group 819:  merge  fork  transition  place  bypass 
    -- CP-element group 819: predecessors 
    -- CP-element group 819: 	808 
    -- CP-element group 819: 	818 
    -- CP-element group 819: successors 
    -- CP-element group 819: 	820 
    -- CP-element group 819: 	821 
    -- CP-element group 819: 	822 
    -- CP-element group 819:  members (2) 
      -- CP-element group 819: 	 branch_block_stmt_714/merge_stmt_1306_PhiReqMerge
      -- CP-element group 819: 	 branch_block_stmt_714/merge_stmt_1306_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(819) <= OrReduce(zeropad3D_CP_2152_elements(808) & zeropad3D_CP_2152_elements(818));
    -- CP-element group 820:  transition  input  bypass 
    -- CP-element group 820: predecessors 
    -- CP-element group 820: 	819 
    -- CP-element group 820: successors 
    -- CP-element group 820: 	823 
    -- CP-element group 820:  members (1) 
      -- CP-element group 820: 	 branch_block_stmt_714/merge_stmt_1306_PhiAck/phi_stmt_1307_ack
      -- 
    phi_stmt_1307_ack_11311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 820_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1307_ack_0, ack => zeropad3D_CP_2152_elements(820)); -- 
    -- CP-element group 821:  transition  input  bypass 
    -- CP-element group 821: predecessors 
    -- CP-element group 821: 	819 
    -- CP-element group 821: successors 
    -- CP-element group 821: 	823 
    -- CP-element group 821:  members (1) 
      -- CP-element group 821: 	 branch_block_stmt_714/merge_stmt_1306_PhiAck/phi_stmt_1313_ack
      -- 
    phi_stmt_1313_ack_11312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 821_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1313_ack_0, ack => zeropad3D_CP_2152_elements(821)); -- 
    -- CP-element group 822:  transition  input  bypass 
    -- CP-element group 822: predecessors 
    -- CP-element group 822: 	819 
    -- CP-element group 822: successors 
    -- CP-element group 822: 	823 
    -- CP-element group 822:  members (1) 
      -- CP-element group 822: 	 branch_block_stmt_714/merge_stmt_1306_PhiAck/phi_stmt_1319_ack
      -- 
    phi_stmt_1319_ack_11313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 822_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1319_ack_0, ack => zeropad3D_CP_2152_elements(822)); -- 
    -- CP-element group 823:  join  transition  bypass 
    -- CP-element group 823: predecessors 
    -- CP-element group 823: 	820 
    -- CP-element group 823: 	821 
    -- CP-element group 823: 	822 
    -- CP-element group 823: successors 
    -- CP-element group 823: 	1 
    -- CP-element group 823:  members (1) 
      -- CP-element group 823: 	 branch_block_stmt_714/merge_stmt_1306_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_823: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_823"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(820) & zeropad3D_CP_2152_elements(821) & zeropad3D_CP_2152_elements(822);
      gj_zeropad3D_cp_element_group_823 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(823), clk => clk, reset => reset); --
    end block;
    -- CP-element group 824:  transition  input  bypass 
    -- CP-element group 824: predecessors 
    -- CP-element group 824: 	133 
    -- CP-element group 824: successors 
    -- CP-element group 824: 	826 
    -- CP-element group 824:  members (2) 
      -- CP-element group 824: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/type_cast_1332/SplitProtocol/Sample/$exit
      -- CP-element group 824: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/type_cast_1332/SplitProtocol/Sample/ra
      -- 
    ra_11333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 824_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1332_inst_ack_0, ack => zeropad3D_CP_2152_elements(824)); -- 
    -- CP-element group 825:  transition  input  bypass 
    -- CP-element group 825: predecessors 
    -- CP-element group 825: 	133 
    -- CP-element group 825: successors 
    -- CP-element group 825: 	826 
    -- CP-element group 825:  members (2) 
      -- CP-element group 825: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/type_cast_1332/SplitProtocol/Update/$exit
      -- CP-element group 825: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/type_cast_1332/SplitProtocol/Update/ca
      -- 
    ca_11338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 825_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1332_inst_ack_1, ack => zeropad3D_CP_2152_elements(825)); -- 
    -- CP-element group 826:  join  transition  output  bypass 
    -- CP-element group 826: predecessors 
    -- CP-element group 826: 	824 
    -- CP-element group 826: 	825 
    -- CP-element group 826: successors 
    -- CP-element group 826: 	830 
    -- CP-element group 826:  members (5) 
      -- CP-element group 826: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/$exit
      -- CP-element group 826: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/$exit
      -- CP-element group 826: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/type_cast_1332/$exit
      -- CP-element group 826: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_sources/type_cast_1332/SplitProtocol/$exit
      -- CP-element group 826: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1329/phi_stmt_1329_req
      -- 
    phi_stmt_1329_req_11339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1329_req_11339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(826), ack => phi_stmt_1329_req_0); -- 
    zeropad3D_cp_element_group_826: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_826"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(824) & zeropad3D_CP_2152_elements(825);
      gj_zeropad3D_cp_element_group_826 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(826), clk => clk, reset => reset); --
    end block;
    -- CP-element group 827:  transition  input  bypass 
    -- CP-element group 827: predecessors 
    -- CP-element group 827: 	133 
    -- CP-element group 827: successors 
    -- CP-element group 827: 	829 
    -- CP-element group 827:  members (2) 
      -- CP-element group 827: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/type_cast_1336/SplitProtocol/Sample/$exit
      -- CP-element group 827: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/type_cast_1336/SplitProtocol/Sample/ra
      -- 
    ra_11356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 827_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1336_inst_ack_0, ack => zeropad3D_CP_2152_elements(827)); -- 
    -- CP-element group 828:  transition  input  bypass 
    -- CP-element group 828: predecessors 
    -- CP-element group 828: 	133 
    -- CP-element group 828: successors 
    -- CP-element group 828: 	829 
    -- CP-element group 828:  members (2) 
      -- CP-element group 828: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/type_cast_1336/SplitProtocol/Update/$exit
      -- CP-element group 828: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/type_cast_1336/SplitProtocol/Update/ca
      -- 
    ca_11361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 828_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1336_inst_ack_1, ack => zeropad3D_CP_2152_elements(828)); -- 
    -- CP-element group 829:  join  transition  output  bypass 
    -- CP-element group 829: predecessors 
    -- CP-element group 829: 	827 
    -- CP-element group 829: 	828 
    -- CP-element group 829: successors 
    -- CP-element group 829: 	830 
    -- CP-element group 829:  members (5) 
      -- CP-element group 829: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/$exit
      -- CP-element group 829: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/$exit
      -- CP-element group 829: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/type_cast_1336/$exit
      -- CP-element group 829: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_sources/type_cast_1336/SplitProtocol/$exit
      -- CP-element group 829: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/phi_stmt_1333/phi_stmt_1333_req
      -- 
    phi_stmt_1333_req_11362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1333_req_11362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(829), ack => phi_stmt_1333_req_0); -- 
    zeropad3D_cp_element_group_829: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_829"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(827) & zeropad3D_CP_2152_elements(828);
      gj_zeropad3D_cp_element_group_829 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(829), clk => clk, reset => reset); --
    end block;
    -- CP-element group 830:  join  fork  transition  place  bypass 
    -- CP-element group 830: predecessors 
    -- CP-element group 830: 	826 
    -- CP-element group 830: 	829 
    -- CP-element group 830: successors 
    -- CP-element group 830: 	831 
    -- CP-element group 830: 	832 
    -- CP-element group 830:  members (3) 
      -- CP-element group 830: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/$exit
      -- CP-element group 830: 	 branch_block_stmt_714/merge_stmt_1328_PhiReqMerge
      -- CP-element group 830: 	 branch_block_stmt_714/merge_stmt_1328_PhiAck/$entry
      -- 
    zeropad3D_cp_element_group_830: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_830"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(826) & zeropad3D_CP_2152_elements(829);
      gj_zeropad3D_cp_element_group_830 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(830), clk => clk, reset => reset); --
    end block;
    -- CP-element group 831:  transition  input  bypass 
    -- CP-element group 831: predecessors 
    -- CP-element group 831: 	830 
    -- CP-element group 831: successors 
    -- CP-element group 831: 	833 
    -- CP-element group 831:  members (1) 
      -- CP-element group 831: 	 branch_block_stmt_714/merge_stmt_1328_PhiAck/phi_stmt_1329_ack
      -- 
    phi_stmt_1329_ack_11367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 831_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1329_ack_0, ack => zeropad3D_CP_2152_elements(831)); -- 
    -- CP-element group 832:  transition  input  bypass 
    -- CP-element group 832: predecessors 
    -- CP-element group 832: 	830 
    -- CP-element group 832: successors 
    -- CP-element group 832: 	833 
    -- CP-element group 832:  members (1) 
      -- CP-element group 832: 	 branch_block_stmt_714/merge_stmt_1328_PhiAck/phi_stmt_1333_ack
      -- 
    phi_stmt_1333_ack_11368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 832_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1333_ack_0, ack => zeropad3D_CP_2152_elements(832)); -- 
    -- CP-element group 833:  join  fork  transition  place  output  bypass 
    -- CP-element group 833: predecessors 
    -- CP-element group 833: 	831 
    -- CP-element group 833: 	832 
    -- CP-element group 833: successors 
    -- CP-element group 833: 	135 
    -- CP-element group 833: 	136 
    -- CP-element group 833: 	137 
    -- CP-element group 833: 	138 
    -- CP-element group 833: 	139 
    -- CP-element group 833: 	140 
    -- CP-element group 833: 	141 
    -- CP-element group 833: 	142 
    -- CP-element group 833: 	143 
    -- CP-element group 833: 	144 
    -- CP-element group 833: 	146 
    -- CP-element group 833: 	148 
    -- CP-element group 833:  members (92) 
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461__entry__
      -- CP-element group 833: 	 branch_block_stmt_714/merge_stmt_1328__exit__
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1340_sample_start_
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1340_update_start_
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1340_Sample/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1340_Sample/rr
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1340_Update/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1340_Update/cr
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_sample_start_
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_update_start_
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_word_address_calculated
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_root_address_calculated
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Sample/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Sample/word_access_start/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Sample/word_access_start/word_0/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Sample/word_access_start/word_0/rr
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Update/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Update/word_access_complete/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Update/word_access_complete/word_0/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_pad_1349_Update/word_access_complete/word_0/cr
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_sample_start_
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_update_start_
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_word_address_calculated
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_root_address_calculated
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Sample/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Sample/word_access_start/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Sample/word_access_start/word_0/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Sample/word_access_start/word_0/rr
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Update/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Update/word_access_complete/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Update/word_access_complete/word_0/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/LOAD_depth_high_1352_Update/word_access_complete/word_0/cr
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_sample_start_
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_update_start_
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_base_address_calculated
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_word_address_calculated
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_root_address_calculated
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_base_address_resized
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_base_addr_resize/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_base_addr_resize/$exit
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_base_addr_resize/base_resize_req
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_base_addr_resize/base_resize_ack
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_base_plus_offset/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_base_plus_offset/$exit
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_base_plus_offset/sum_rename_req
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_base_plus_offset/sum_rename_ack
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_word_addrgen/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_word_addrgen/$exit
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_word_addrgen/root_register_req
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_word_addrgen/root_register_ack
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Sample/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Sample/word_access_start/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Sample/word_access_start/word_0/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Sample/word_access_start/word_0/rr
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Update/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Update/word_access_complete/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Update/word_access_complete/word_0/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1364_Update/word_access_complete/word_0/cr
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_sample_start_
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_update_start_
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_base_address_calculated
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_word_address_calculated
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_root_address_calculated
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_base_address_resized
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_base_addr_resize/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_base_addr_resize/$exit
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_base_addr_resize/base_resize_req
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_base_addr_resize/base_resize_ack
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_base_plus_offset/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_base_plus_offset/$exit
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_base_plus_offset/sum_rename_req
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_base_plus_offset/sum_rename_ack
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_word_addrgen/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_word_addrgen/$exit
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_word_addrgen/root_register_req
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_word_addrgen/root_register_ack
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Sample/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Sample/word_access_start/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Sample/word_access_start/word_0/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Sample/word_access_start/word_0/rr
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Update/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Update/word_access_complete/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Update/word_access_complete/word_0/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/ptr_deref_1376_Update/word_access_complete/word_0/cr
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1380_update_start_
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1380_Update/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1380_Update/cr
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1419_update_start_
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1419_Update/$entry
      -- CP-element group 833: 	 branch_block_stmt_714/assign_stmt_1341_to_assign_stmt_1461/type_cast_1419_Update/cr
      -- CP-element group 833: 	 branch_block_stmt_714/merge_stmt_1328_PhiAck/$exit
      -- 
    rr_3951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(833), ack => type_cast_1340_inst_req_0); -- 
    cr_3956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(833), ack => type_cast_1340_inst_req_1); -- 
    rr_3973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(833), ack => LOAD_pad_1349_load_0_req_0); -- 
    cr_3984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(833), ack => LOAD_pad_1349_load_0_req_1); -- 
    rr_4006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(833), ack => LOAD_depth_high_1352_load_0_req_0); -- 
    cr_4017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(833), ack => LOAD_depth_high_1352_load_0_req_1); -- 
    rr_4056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(833), ack => ptr_deref_1364_load_0_req_0); -- 
    cr_4067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(833), ack => ptr_deref_1364_load_0_req_1); -- 
    rr_4106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(833), ack => ptr_deref_1376_load_0_req_0); -- 
    cr_4117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(833), ack => ptr_deref_1376_load_0_req_1); -- 
    cr_4136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(833), ack => type_cast_1380_inst_req_1); -- 
    cr_4150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(833), ack => type_cast_1419_inst_req_1); -- 
    zeropad3D_cp_element_group_833: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_833"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(831) & zeropad3D_CP_2152_elements(832);
      gj_zeropad3D_cp_element_group_833 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(833), clk => clk, reset => reset); --
    end block;
    -- CP-element group 834:  transition  input  bypass 
    -- CP-element group 834: predecessors 
    -- CP-element group 834: 	2 
    -- CP-element group 834: successors 
    -- CP-element group 834: 	836 
    -- CP-element group 834:  members (2) 
      -- CP-element group 834: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1469/SplitProtocol/Sample/$exit
      -- CP-element group 834: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1469/SplitProtocol/Sample/ra
      -- 
    ra_11388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 834_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1469_inst_ack_0, ack => zeropad3D_CP_2152_elements(834)); -- 
    -- CP-element group 835:  transition  input  bypass 
    -- CP-element group 835: predecessors 
    -- CP-element group 835: 	2 
    -- CP-element group 835: successors 
    -- CP-element group 835: 	836 
    -- CP-element group 835:  members (2) 
      -- CP-element group 835: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1469/SplitProtocol/Update/$exit
      -- CP-element group 835: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1469/SplitProtocol/Update/ca
      -- 
    ca_11393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 835_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1469_inst_ack_1, ack => zeropad3D_CP_2152_elements(835)); -- 
    -- CP-element group 836:  join  transition  output  bypass 
    -- CP-element group 836: predecessors 
    -- CP-element group 836: 	834 
    -- CP-element group 836: 	835 
    -- CP-element group 836: successors 
    -- CP-element group 836: 	843 
    -- CP-element group 836:  members (5) 
      -- CP-element group 836: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/$exit
      -- CP-element group 836: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/$exit
      -- CP-element group 836: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1469/$exit
      -- CP-element group 836: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1469/SplitProtocol/$exit
      -- CP-element group 836: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_req
      -- 
    phi_stmt_1464_req_11394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1464_req_11394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(836), ack => phi_stmt_1464_req_1); -- 
    zeropad3D_cp_element_group_836: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_836"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(834) & zeropad3D_CP_2152_elements(835);
      gj_zeropad3D_cp_element_group_836 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(836), clk => clk, reset => reset); --
    end block;
    -- CP-element group 837:  transition  input  bypass 
    -- CP-element group 837: predecessors 
    -- CP-element group 837: 	2 
    -- CP-element group 837: successors 
    -- CP-element group 837: 	839 
    -- CP-element group 837:  members (2) 
      -- CP-element group 837: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/type_cast_1476/SplitProtocol/Sample/$exit
      -- CP-element group 837: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/type_cast_1476/SplitProtocol/Sample/ra
      -- 
    ra_11411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 837_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1476_inst_ack_0, ack => zeropad3D_CP_2152_elements(837)); -- 
    -- CP-element group 838:  transition  input  bypass 
    -- CP-element group 838: predecessors 
    -- CP-element group 838: 	2 
    -- CP-element group 838: successors 
    -- CP-element group 838: 	839 
    -- CP-element group 838:  members (2) 
      -- CP-element group 838: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/type_cast_1476/SplitProtocol/Update/$exit
      -- CP-element group 838: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/type_cast_1476/SplitProtocol/Update/ca
      -- 
    ca_11416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 838_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1476_inst_ack_1, ack => zeropad3D_CP_2152_elements(838)); -- 
    -- CP-element group 839:  join  transition  output  bypass 
    -- CP-element group 839: predecessors 
    -- CP-element group 839: 	837 
    -- CP-element group 839: 	838 
    -- CP-element group 839: successors 
    -- CP-element group 839: 	843 
    -- CP-element group 839:  members (5) 
      -- CP-element group 839: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/$exit
      -- CP-element group 839: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/$exit
      -- CP-element group 839: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/type_cast_1476/$exit
      -- CP-element group 839: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/type_cast_1476/SplitProtocol/$exit
      -- CP-element group 839: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_req
      -- 
    phi_stmt_1470_req_11417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1470_req_11417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(839), ack => phi_stmt_1470_req_1); -- 
    zeropad3D_cp_element_group_839: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_839"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(837) & zeropad3D_CP_2152_elements(838);
      gj_zeropad3D_cp_element_group_839 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(839), clk => clk, reset => reset); --
    end block;
    -- CP-element group 840:  transition  input  bypass 
    -- CP-element group 840: predecessors 
    -- CP-element group 840: 	2 
    -- CP-element group 840: successors 
    -- CP-element group 840: 	842 
    -- CP-element group 840:  members (2) 
      -- CP-element group 840: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/type_cast_1483/SplitProtocol/Sample/$exit
      -- CP-element group 840: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/type_cast_1483/SplitProtocol/Sample/ra
      -- 
    ra_11434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 840_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1483_inst_ack_0, ack => zeropad3D_CP_2152_elements(840)); -- 
    -- CP-element group 841:  transition  input  bypass 
    -- CP-element group 841: predecessors 
    -- CP-element group 841: 	2 
    -- CP-element group 841: successors 
    -- CP-element group 841: 	842 
    -- CP-element group 841:  members (2) 
      -- CP-element group 841: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/type_cast_1483/SplitProtocol/Update/$exit
      -- CP-element group 841: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/type_cast_1483/SplitProtocol/Update/ca
      -- 
    ca_11439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 841_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1483_inst_ack_1, ack => zeropad3D_CP_2152_elements(841)); -- 
    -- CP-element group 842:  join  transition  output  bypass 
    -- CP-element group 842: predecessors 
    -- CP-element group 842: 	840 
    -- CP-element group 842: 	841 
    -- CP-element group 842: successors 
    -- CP-element group 842: 	843 
    -- CP-element group 842:  members (5) 
      -- CP-element group 842: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/$exit
      -- CP-element group 842: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/$exit
      -- CP-element group 842: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/type_cast_1483/$exit
      -- CP-element group 842: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/type_cast_1483/SplitProtocol/$exit
      -- CP-element group 842: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_req
      -- 
    phi_stmt_1477_req_11440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1477_req_11440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(842), ack => phi_stmt_1477_req_1); -- 
    zeropad3D_cp_element_group_842: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_842"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(840) & zeropad3D_CP_2152_elements(841);
      gj_zeropad3D_cp_element_group_842 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(842), clk => clk, reset => reset); --
    end block;
    -- CP-element group 843:  join  transition  bypass 
    -- CP-element group 843: predecessors 
    -- CP-element group 843: 	836 
    -- CP-element group 843: 	839 
    -- CP-element group 843: 	842 
    -- CP-element group 843: successors 
    -- CP-element group 843: 	850 
    -- CP-element group 843:  members (1) 
      -- CP-element group 843: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_843: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_843"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(836) & zeropad3D_CP_2152_elements(839) & zeropad3D_CP_2152_elements(842);
      gj_zeropad3D_cp_element_group_843 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(843), clk => clk, reset => reset); --
    end block;
    -- CP-element group 844:  transition  input  bypass 
    -- CP-element group 844: predecessors 
    -- CP-element group 844: 	149 
    -- CP-element group 844: successors 
    -- CP-element group 844: 	846 
    -- CP-element group 844:  members (2) 
      -- CP-element group 844: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Sample/$exit
      -- CP-element group 844: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Sample/ra
      -- 
    ra_11460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 844_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1467_inst_ack_0, ack => zeropad3D_CP_2152_elements(844)); -- 
    -- CP-element group 845:  transition  input  bypass 
    -- CP-element group 845: predecessors 
    -- CP-element group 845: 	149 
    -- CP-element group 845: successors 
    -- CP-element group 845: 	846 
    -- CP-element group 845:  members (2) 
      -- CP-element group 845: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Update/$exit
      -- CP-element group 845: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/Update/ca
      -- 
    ca_11465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 845_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1467_inst_ack_1, ack => zeropad3D_CP_2152_elements(845)); -- 
    -- CP-element group 846:  join  transition  output  bypass 
    -- CP-element group 846: predecessors 
    -- CP-element group 846: 	844 
    -- CP-element group 846: 	845 
    -- CP-element group 846: successors 
    -- CP-element group 846: 	849 
    -- CP-element group 846:  members (5) 
      -- CP-element group 846: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/$exit
      -- CP-element group 846: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/$exit
      -- CP-element group 846: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/$exit
      -- CP-element group 846: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_sources/type_cast_1467/SplitProtocol/$exit
      -- CP-element group 846: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1464/phi_stmt_1464_req
      -- 
    phi_stmt_1464_req_11466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1464_req_11466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(846), ack => phi_stmt_1464_req_0); -- 
    zeropad3D_cp_element_group_846: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_846"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(844) & zeropad3D_CP_2152_elements(845);
      gj_zeropad3D_cp_element_group_846 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(846), clk => clk, reset => reset); --
    end block;
    -- CP-element group 847:  transition  output  delay-element  bypass 
    -- CP-element group 847: predecessors 
    -- CP-element group 847: 	149 
    -- CP-element group 847: successors 
    -- CP-element group 847: 	849 
    -- CP-element group 847:  members (4) 
      -- CP-element group 847: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1470/$exit
      -- CP-element group 847: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/$exit
      -- CP-element group 847: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_sources/type_cast_1474_konst_delay_trans
      -- CP-element group 847: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1470/phi_stmt_1470_req
      -- 
    phi_stmt_1470_req_11474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1470_req_11474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(847), ack => phi_stmt_1470_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(847) is a control-delay.
    cp_element_847_delay: control_delay_element  generic map(name => " 847_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(149), ack => zeropad3D_CP_2152_elements(847), clk => clk, reset =>reset);
    -- CP-element group 848:  transition  output  delay-element  bypass 
    -- CP-element group 848: predecessors 
    -- CP-element group 848: 	149 
    -- CP-element group 848: successors 
    -- CP-element group 848: 	849 
    -- CP-element group 848:  members (4) 
      -- CP-element group 848: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1477/$exit
      -- CP-element group 848: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/$exit
      -- CP-element group 848: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_sources/type_cast_1481_konst_delay_trans
      -- CP-element group 848: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1477/phi_stmt_1477_req
      -- 
    phi_stmt_1477_req_11482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1477_req_11482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(848), ack => phi_stmt_1477_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(848) is a control-delay.
    cp_element_848_delay: control_delay_element  generic map(name => " 848_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(149), ack => zeropad3D_CP_2152_elements(848), clk => clk, reset =>reset);
    -- CP-element group 849:  join  transition  bypass 
    -- CP-element group 849: predecessors 
    -- CP-element group 849: 	846 
    -- CP-element group 849: 	847 
    -- CP-element group 849: 	848 
    -- CP-element group 849: successors 
    -- CP-element group 849: 	850 
    -- CP-element group 849:  members (1) 
      -- CP-element group 849: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_849: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_849"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(846) & zeropad3D_CP_2152_elements(847) & zeropad3D_CP_2152_elements(848);
      gj_zeropad3D_cp_element_group_849 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(849), clk => clk, reset => reset); --
    end block;
    -- CP-element group 850:  merge  fork  transition  place  bypass 
    -- CP-element group 850: predecessors 
    -- CP-element group 850: 	843 
    -- CP-element group 850: 	849 
    -- CP-element group 850: successors 
    -- CP-element group 850: 	851 
    -- CP-element group 850: 	852 
    -- CP-element group 850: 	853 
    -- CP-element group 850:  members (2) 
      -- CP-element group 850: 	 branch_block_stmt_714/merge_stmt_1463_PhiReqMerge
      -- CP-element group 850: 	 branch_block_stmt_714/merge_stmt_1463_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(850) <= OrReduce(zeropad3D_CP_2152_elements(843) & zeropad3D_CP_2152_elements(849));
    -- CP-element group 851:  transition  input  bypass 
    -- CP-element group 851: predecessors 
    -- CP-element group 851: 	850 
    -- CP-element group 851: successors 
    -- CP-element group 851: 	854 
    -- CP-element group 851:  members (1) 
      -- CP-element group 851: 	 branch_block_stmt_714/merge_stmt_1463_PhiAck/phi_stmt_1464_ack
      -- 
    phi_stmt_1464_ack_11487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 851_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1464_ack_0, ack => zeropad3D_CP_2152_elements(851)); -- 
    -- CP-element group 852:  transition  input  bypass 
    -- CP-element group 852: predecessors 
    -- CP-element group 852: 	850 
    -- CP-element group 852: successors 
    -- CP-element group 852: 	854 
    -- CP-element group 852:  members (1) 
      -- CP-element group 852: 	 branch_block_stmt_714/merge_stmt_1463_PhiAck/phi_stmt_1470_ack
      -- 
    phi_stmt_1470_ack_11488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 852_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1470_ack_0, ack => zeropad3D_CP_2152_elements(852)); -- 
    -- CP-element group 853:  transition  input  bypass 
    -- CP-element group 853: predecessors 
    -- CP-element group 853: 	850 
    -- CP-element group 853: successors 
    -- CP-element group 853: 	854 
    -- CP-element group 853:  members (1) 
      -- CP-element group 853: 	 branch_block_stmt_714/merge_stmt_1463_PhiAck/phi_stmt_1477_ack
      -- 
    phi_stmt_1477_ack_11489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 853_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1477_ack_0, ack => zeropad3D_CP_2152_elements(853)); -- 
    -- CP-element group 854:  join  fork  transition  place  output  bypass 
    -- CP-element group 854: predecessors 
    -- CP-element group 854: 	851 
    -- CP-element group 854: 	852 
    -- CP-element group 854: 	853 
    -- CP-element group 854: successors 
    -- CP-element group 854: 	150 
    -- CP-element group 854: 	151 
    -- CP-element group 854:  members (10) 
      -- CP-element group 854: 	 branch_block_stmt_714/merge_stmt_1463__exit__
      -- CP-element group 854: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496__entry__
      -- CP-element group 854: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/$entry
      -- CP-element group 854: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/type_cast_1488_sample_start_
      -- CP-element group 854: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/type_cast_1488_update_start_
      -- CP-element group 854: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/type_cast_1488_Sample/$entry
      -- CP-element group 854: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/type_cast_1488_Sample/rr
      -- CP-element group 854: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/type_cast_1488_Update/$entry
      -- CP-element group 854: 	 branch_block_stmt_714/assign_stmt_1489_to_assign_stmt_1496/type_cast_1488_Update/cr
      -- CP-element group 854: 	 branch_block_stmt_714/merge_stmt_1463_PhiAck/$exit
      -- 
    rr_4162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(854), ack => type_cast_1488_inst_req_0); -- 
    cr_4167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(854), ack => type_cast_1488_inst_req_1); -- 
    zeropad3D_cp_element_group_854: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_854"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(851) & zeropad3D_CP_2152_elements(852) & zeropad3D_CP_2152_elements(853);
      gj_zeropad3D_cp_element_group_854 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(854), clk => clk, reset => reset); --
    end block;
    -- CP-element group 855:  merge  fork  transition  place  output  bypass 
    -- CP-element group 855: predecessors 
    -- CP-element group 855: 	152 
    -- CP-element group 855: 	159 
    -- CP-element group 855: 	162 
    -- CP-element group 855: 	169 
    -- CP-element group 855: successors 
    -- CP-element group 855: 	170 
    -- CP-element group 855: 	171 
    -- CP-element group 855: 	172 
    -- CP-element group 855: 	173 
    -- CP-element group 855: 	176 
    -- CP-element group 855: 	178 
    -- CP-element group 855: 	180 
    -- CP-element group 855: 	182 
    -- CP-element group 855:  members (33) 
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636__entry__
      -- CP-element group 855: 	 branch_block_stmt_714/merge_stmt_1580__exit__
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_final_index_sum_regn_update_start
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/$entry
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/addr_of_1630_update_start_
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1623_Update/cr
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_update_start_
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Update/word_access_complete/word_0/cr
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1623_Update/$entry
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/addr_of_1630_complete/req
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Update/word_access_complete/word_0/$entry
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Update/word_access_complete/$entry
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/addr_of_1630_complete/$entry
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1623_update_start_
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1589_Update/cr
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/ptr_deref_1633_Update/$entry
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1589_Update/$entry
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1589_Sample/rr
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1589_Sample/$entry
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1589_update_start_
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1589_sample_start_
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1584_Update/cr
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1584_Update/$entry
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1584_Sample/rr
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_final_index_sum_regn_Update/req
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/array_obj_ref_1629_final_index_sum_regn_Update/$entry
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1584_Sample/$entry
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1584_update_start_
      -- CP-element group 855: 	 branch_block_stmt_714/assign_stmt_1585_to_assign_stmt_1636/type_cast_1584_sample_start_
      -- CP-element group 855: 	 branch_block_stmt_714/merge_stmt_1580_PhiReqMerge
      -- CP-element group 855: 	 branch_block_stmt_714/merge_stmt_1580_PhiAck/$entry
      -- CP-element group 855: 	 branch_block_stmt_714/merge_stmt_1580_PhiAck/$exit
      -- CP-element group 855: 	 branch_block_stmt_714/merge_stmt_1580_PhiAck/dummy
      -- 
    cr_4405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(855), ack => type_cast_1623_inst_req_1); -- 
    cr_4501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(855), ack => ptr_deref_1633_store_0_req_1); -- 
    req_4451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(855), ack => addr_of_1630_final_reg_req_1); -- 
    cr_4391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(855), ack => type_cast_1589_inst_req_1); -- 
    rr_4386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(855), ack => type_cast_1589_inst_req_0); -- 
    cr_4377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(855), ack => type_cast_1584_inst_req_1); -- 
    rr_4372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(855), ack => type_cast_1584_inst_req_0); -- 
    req_4436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(855), ack => array_obj_ref_1629_index_offset_req_1); -- 
    zeropad3D_CP_2152_elements(855) <= OrReduce(zeropad3D_CP_2152_elements(152) & zeropad3D_CP_2152_elements(159) & zeropad3D_CP_2152_elements(162) & zeropad3D_CP_2152_elements(169));
    -- CP-element group 856:  merge  fork  transition  place  output  bypass 
    -- CP-element group 856: predecessors 
    -- CP-element group 856: 	183 
    -- CP-element group 856: 	203 
    -- CP-element group 856: successors 
    -- CP-element group 856: 	204 
    -- CP-element group 856: 	205 
    -- CP-element group 856:  members (13) 
      -- CP-element group 856: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763__entry__
      -- CP-element group 856: 	 branch_block_stmt_714/merge_stmt_1745__exit__
      -- CP-element group 856: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/$entry
      -- CP-element group 856: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/type_cast_1749_sample_start_
      -- CP-element group 856: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/type_cast_1749_update_start_
      -- CP-element group 856: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/type_cast_1749_Sample/$entry
      -- CP-element group 856: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/type_cast_1749_Sample/rr
      -- CP-element group 856: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/type_cast_1749_Update/$entry
      -- CP-element group 856: 	 branch_block_stmt_714/assign_stmt_1750_to_assign_stmt_1763/type_cast_1749_Update/cr
      -- CP-element group 856: 	 branch_block_stmt_714/merge_stmt_1745_PhiReqMerge
      -- CP-element group 856: 	 branch_block_stmt_714/merge_stmt_1745_PhiAck/$entry
      -- CP-element group 856: 	 branch_block_stmt_714/merge_stmt_1745_PhiAck/$exit
      -- CP-element group 856: 	 branch_block_stmt_714/merge_stmt_1745_PhiAck/dummy
      -- 
    rr_4750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(856), ack => type_cast_1749_inst_req_0); -- 
    cr_4755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(856), ack => type_cast_1749_inst_req_1); -- 
    zeropad3D_CP_2152_elements(856) <= OrReduce(zeropad3D_CP_2152_elements(183) & zeropad3D_CP_2152_elements(203));
    -- CP-element group 857:  transition  output  delay-element  bypass 
    -- CP-element group 857: predecessors 
    -- CP-element group 857: 	225 
    -- CP-element group 857: successors 
    -- CP-element group 857: 	864 
    -- CP-element group 857:  members (4) 
      -- CP-element group 857: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1869/$exit
      -- CP-element group 857: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/$exit
      -- CP-element group 857: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/type_cast_1875_konst_delay_trans
      -- CP-element group 857: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_req
      -- 
    phi_stmt_1869_req_11600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1869_req_11600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(857), ack => phi_stmt_1869_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(857) is a control-delay.
    cp_element_857_delay: control_delay_element  generic map(name => " 857_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(225), ack => zeropad3D_CP_2152_elements(857), clk => clk, reset =>reset);
    -- CP-element group 858:  transition  input  bypass 
    -- CP-element group 858: predecessors 
    -- CP-element group 858: 	225 
    -- CP-element group 858: successors 
    -- CP-element group 858: 	860 
    -- CP-element group 858:  members (2) 
      -- CP-element group 858: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1868/SplitProtocol/Sample/$exit
      -- CP-element group 858: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1868/SplitProtocol/Sample/ra
      -- 
    ra_11617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 858_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1868_inst_ack_0, ack => zeropad3D_CP_2152_elements(858)); -- 
    -- CP-element group 859:  transition  input  bypass 
    -- CP-element group 859: predecessors 
    -- CP-element group 859: 	225 
    -- CP-element group 859: successors 
    -- CP-element group 859: 	860 
    -- CP-element group 859:  members (2) 
      -- CP-element group 859: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1868/SplitProtocol/Update/$exit
      -- CP-element group 859: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1868/SplitProtocol/Update/ca
      -- 
    ca_11622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 859_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1868_inst_ack_1, ack => zeropad3D_CP_2152_elements(859)); -- 
    -- CP-element group 860:  join  transition  output  bypass 
    -- CP-element group 860: predecessors 
    -- CP-element group 860: 	858 
    -- CP-element group 860: 	859 
    -- CP-element group 860: successors 
    -- CP-element group 860: 	864 
    -- CP-element group 860:  members (5) 
      -- CP-element group 860: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/$exit
      -- CP-element group 860: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/$exit
      -- CP-element group 860: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1868/$exit
      -- CP-element group 860: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1868/SplitProtocol/$exit
      -- CP-element group 860: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_req
      -- 
    phi_stmt_1863_req_11623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1863_req_11623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(860), ack => phi_stmt_1863_req_1); -- 
    zeropad3D_cp_element_group_860: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_860"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(858) & zeropad3D_CP_2152_elements(859);
      gj_zeropad3D_cp_element_group_860 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(860), clk => clk, reset => reset); --
    end block;
    -- CP-element group 861:  transition  input  bypass 
    -- CP-element group 861: predecessors 
    -- CP-element group 861: 	225 
    -- CP-element group 861: successors 
    -- CP-element group 861: 	863 
    -- CP-element group 861:  members (2) 
      -- CP-element group 861: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1862/SplitProtocol/Sample/$exit
      -- CP-element group 861: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1862/SplitProtocol/Sample/ra
      -- 
    ra_11640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 861_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1862_inst_ack_0, ack => zeropad3D_CP_2152_elements(861)); -- 
    -- CP-element group 862:  transition  input  bypass 
    -- CP-element group 862: predecessors 
    -- CP-element group 862: 	225 
    -- CP-element group 862: successors 
    -- CP-element group 862: 	863 
    -- CP-element group 862:  members (2) 
      -- CP-element group 862: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1862/SplitProtocol/Update/$exit
      -- CP-element group 862: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1862/SplitProtocol/Update/ca
      -- 
    ca_11645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 862_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1862_inst_ack_1, ack => zeropad3D_CP_2152_elements(862)); -- 
    -- CP-element group 863:  join  transition  output  bypass 
    -- CP-element group 863: predecessors 
    -- CP-element group 863: 	861 
    -- CP-element group 863: 	862 
    -- CP-element group 863: successors 
    -- CP-element group 863: 	864 
    -- CP-element group 863:  members (5) 
      -- CP-element group 863: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/$exit
      -- CP-element group 863: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/$exit
      -- CP-element group 863: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1862/$exit
      -- CP-element group 863: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1862/SplitProtocol/$exit
      -- CP-element group 863: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_req
      -- 
    phi_stmt_1857_req_11646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1857_req_11646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(863), ack => phi_stmt_1857_req_1); -- 
    zeropad3D_cp_element_group_863: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_863"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(861) & zeropad3D_CP_2152_elements(862);
      gj_zeropad3D_cp_element_group_863 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(863), clk => clk, reset => reset); --
    end block;
    -- CP-element group 864:  join  transition  bypass 
    -- CP-element group 864: predecessors 
    -- CP-element group 864: 	857 
    -- CP-element group 864: 	860 
    -- CP-element group 864: 	863 
    -- CP-element group 864: successors 
    -- CP-element group 864: 	875 
    -- CP-element group 864:  members (1) 
      -- CP-element group 864: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_864: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_864"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(857) & zeropad3D_CP_2152_elements(860) & zeropad3D_CP_2152_elements(863);
      gj_zeropad3D_cp_element_group_864 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(864), clk => clk, reset => reset); --
    end block;
    -- CP-element group 865:  transition  input  bypass 
    -- CP-element group 865: predecessors 
    -- CP-element group 865: 	206 
    -- CP-element group 865: successors 
    -- CP-element group 865: 	867 
    -- CP-element group 865:  members (2) 
      -- CP-element group 865: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/type_cast_1872/SplitProtocol/Sample/$exit
      -- CP-element group 865: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/type_cast_1872/SplitProtocol/Sample/ra
      -- 
    ra_11666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 865_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1872_inst_ack_0, ack => zeropad3D_CP_2152_elements(865)); -- 
    -- CP-element group 866:  transition  input  bypass 
    -- CP-element group 866: predecessors 
    -- CP-element group 866: 	206 
    -- CP-element group 866: successors 
    -- CP-element group 866: 	867 
    -- CP-element group 866:  members (2) 
      -- CP-element group 866: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/type_cast_1872/SplitProtocol/Update/$exit
      -- CP-element group 866: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/type_cast_1872/SplitProtocol/Update/ca
      -- 
    ca_11671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 866_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1872_inst_ack_1, ack => zeropad3D_CP_2152_elements(866)); -- 
    -- CP-element group 867:  join  transition  output  bypass 
    -- CP-element group 867: predecessors 
    -- CP-element group 867: 	865 
    -- CP-element group 867: 	866 
    -- CP-element group 867: successors 
    -- CP-element group 867: 	874 
    -- CP-element group 867:  members (5) 
      -- CP-element group 867: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/$exit
      -- CP-element group 867: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/$exit
      -- CP-element group 867: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/type_cast_1872/$exit
      -- CP-element group 867: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_sources/type_cast_1872/SplitProtocol/$exit
      -- CP-element group 867: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1869/phi_stmt_1869_req
      -- 
    phi_stmt_1869_req_11672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1869_req_11672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(867), ack => phi_stmt_1869_req_0); -- 
    zeropad3D_cp_element_group_867: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_867"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(865) & zeropad3D_CP_2152_elements(866);
      gj_zeropad3D_cp_element_group_867 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(867), clk => clk, reset => reset); --
    end block;
    -- CP-element group 868:  transition  input  bypass 
    -- CP-element group 868: predecessors 
    -- CP-element group 868: 	206 
    -- CP-element group 868: successors 
    -- CP-element group 868: 	870 
    -- CP-element group 868:  members (2) 
      -- CP-element group 868: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1866/SplitProtocol/Sample/$exit
      -- CP-element group 868: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1866/SplitProtocol/Sample/ra
      -- 
    ra_11689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 868_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1866_inst_ack_0, ack => zeropad3D_CP_2152_elements(868)); -- 
    -- CP-element group 869:  transition  input  bypass 
    -- CP-element group 869: predecessors 
    -- CP-element group 869: 	206 
    -- CP-element group 869: successors 
    -- CP-element group 869: 	870 
    -- CP-element group 869:  members (2) 
      -- CP-element group 869: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1866/SplitProtocol/Update/$exit
      -- CP-element group 869: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1866/SplitProtocol/Update/ca
      -- 
    ca_11694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 869_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1866_inst_ack_1, ack => zeropad3D_CP_2152_elements(869)); -- 
    -- CP-element group 870:  join  transition  output  bypass 
    -- CP-element group 870: predecessors 
    -- CP-element group 870: 	868 
    -- CP-element group 870: 	869 
    -- CP-element group 870: successors 
    -- CP-element group 870: 	874 
    -- CP-element group 870:  members (5) 
      -- CP-element group 870: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/$exit
      -- CP-element group 870: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/$exit
      -- CP-element group 870: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1866/$exit
      -- CP-element group 870: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_sources/type_cast_1866/SplitProtocol/$exit
      -- CP-element group 870: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1863/phi_stmt_1863_req
      -- 
    phi_stmt_1863_req_11695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1863_req_11695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(870), ack => phi_stmt_1863_req_0); -- 
    zeropad3D_cp_element_group_870: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_870"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(868) & zeropad3D_CP_2152_elements(869);
      gj_zeropad3D_cp_element_group_870 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(870), clk => clk, reset => reset); --
    end block;
    -- CP-element group 871:  transition  input  bypass 
    -- CP-element group 871: predecessors 
    -- CP-element group 871: 	206 
    -- CP-element group 871: successors 
    -- CP-element group 871: 	873 
    -- CP-element group 871:  members (2) 
      -- CP-element group 871: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1860/SplitProtocol/Sample/$exit
      -- CP-element group 871: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1860/SplitProtocol/Sample/ra
      -- 
    ra_11712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 871_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1860_inst_ack_0, ack => zeropad3D_CP_2152_elements(871)); -- 
    -- CP-element group 872:  transition  input  bypass 
    -- CP-element group 872: predecessors 
    -- CP-element group 872: 	206 
    -- CP-element group 872: successors 
    -- CP-element group 872: 	873 
    -- CP-element group 872:  members (2) 
      -- CP-element group 872: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1860/SplitProtocol/Update/$exit
      -- CP-element group 872: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1860/SplitProtocol/Update/ca
      -- 
    ca_11717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 872_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1860_inst_ack_1, ack => zeropad3D_CP_2152_elements(872)); -- 
    -- CP-element group 873:  join  transition  output  bypass 
    -- CP-element group 873: predecessors 
    -- CP-element group 873: 	871 
    -- CP-element group 873: 	872 
    -- CP-element group 873: successors 
    -- CP-element group 873: 	874 
    -- CP-element group 873:  members (5) 
      -- CP-element group 873: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/$exit
      -- CP-element group 873: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/$exit
      -- CP-element group 873: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1860/$exit
      -- CP-element group 873: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_sources/type_cast_1860/SplitProtocol/$exit
      -- CP-element group 873: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1857/phi_stmt_1857_req
      -- 
    phi_stmt_1857_req_11718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1857_req_11718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(873), ack => phi_stmt_1857_req_0); -- 
    zeropad3D_cp_element_group_873: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_873"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(871) & zeropad3D_CP_2152_elements(872);
      gj_zeropad3D_cp_element_group_873 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(873), clk => clk, reset => reset); --
    end block;
    -- CP-element group 874:  join  transition  bypass 
    -- CP-element group 874: predecessors 
    -- CP-element group 874: 	867 
    -- CP-element group 874: 	870 
    -- CP-element group 874: 	873 
    -- CP-element group 874: successors 
    -- CP-element group 874: 	875 
    -- CP-element group 874:  members (1) 
      -- CP-element group 874: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_874: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_874"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(867) & zeropad3D_CP_2152_elements(870) & zeropad3D_CP_2152_elements(873);
      gj_zeropad3D_cp_element_group_874 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(874), clk => clk, reset => reset); --
    end block;
    -- CP-element group 875:  merge  fork  transition  place  bypass 
    -- CP-element group 875: predecessors 
    -- CP-element group 875: 	864 
    -- CP-element group 875: 	874 
    -- CP-element group 875: successors 
    -- CP-element group 875: 	876 
    -- CP-element group 875: 	877 
    -- CP-element group 875: 	878 
    -- CP-element group 875:  members (2) 
      -- CP-element group 875: 	 branch_block_stmt_714/merge_stmt_1856_PhiReqMerge
      -- CP-element group 875: 	 branch_block_stmt_714/merge_stmt_1856_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(875) <= OrReduce(zeropad3D_CP_2152_elements(864) & zeropad3D_CP_2152_elements(874));
    -- CP-element group 876:  transition  input  bypass 
    -- CP-element group 876: predecessors 
    -- CP-element group 876: 	875 
    -- CP-element group 876: successors 
    -- CP-element group 876: 	879 
    -- CP-element group 876:  members (1) 
      -- CP-element group 876: 	 branch_block_stmt_714/merge_stmt_1856_PhiAck/phi_stmt_1857_ack
      -- 
    phi_stmt_1857_ack_11723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 876_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1857_ack_0, ack => zeropad3D_CP_2152_elements(876)); -- 
    -- CP-element group 877:  transition  input  bypass 
    -- CP-element group 877: predecessors 
    -- CP-element group 877: 	875 
    -- CP-element group 877: successors 
    -- CP-element group 877: 	879 
    -- CP-element group 877:  members (1) 
      -- CP-element group 877: 	 branch_block_stmt_714/merge_stmt_1856_PhiAck/phi_stmt_1863_ack
      -- 
    phi_stmt_1863_ack_11724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 877_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1863_ack_0, ack => zeropad3D_CP_2152_elements(877)); -- 
    -- CP-element group 878:  transition  input  bypass 
    -- CP-element group 878: predecessors 
    -- CP-element group 878: 	875 
    -- CP-element group 878: successors 
    -- CP-element group 878: 	879 
    -- CP-element group 878:  members (1) 
      -- CP-element group 878: 	 branch_block_stmt_714/merge_stmt_1856_PhiAck/phi_stmt_1869_ack
      -- 
    phi_stmt_1869_ack_11725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 878_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1869_ack_0, ack => zeropad3D_CP_2152_elements(878)); -- 
    -- CP-element group 879:  join  transition  bypass 
    -- CP-element group 879: predecessors 
    -- CP-element group 879: 	876 
    -- CP-element group 879: 	877 
    -- CP-element group 879: 	878 
    -- CP-element group 879: successors 
    -- CP-element group 879: 	2 
    -- CP-element group 879:  members (1) 
      -- CP-element group 879: 	 branch_block_stmt_714/merge_stmt_1856_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_879: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_879"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(876) & zeropad3D_CP_2152_elements(877) & zeropad3D_CP_2152_elements(878);
      gj_zeropad3D_cp_element_group_879 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(879), clk => clk, reset => reset); --
    end block;
    -- CP-element group 880:  transition  input  bypass 
    -- CP-element group 880: predecessors 
    -- CP-element group 880: 	224 
    -- CP-element group 880: successors 
    -- CP-element group 880: 	882 
    -- CP-element group 880:  members (2) 
      -- CP-element group 880: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/type_cast_1886/SplitProtocol/Sample/$exit
      -- CP-element group 880: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/type_cast_1886/SplitProtocol/Sample/ra
      -- 
    ra_11745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 880_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1886_inst_ack_0, ack => zeropad3D_CP_2152_elements(880)); -- 
    -- CP-element group 881:  transition  input  bypass 
    -- CP-element group 881: predecessors 
    -- CP-element group 881: 	224 
    -- CP-element group 881: successors 
    -- CP-element group 881: 	882 
    -- CP-element group 881:  members (2) 
      -- CP-element group 881: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/type_cast_1886/SplitProtocol/Update/$exit
      -- CP-element group 881: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/type_cast_1886/SplitProtocol/Update/ca
      -- 
    ca_11750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 881_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1886_inst_ack_1, ack => zeropad3D_CP_2152_elements(881)); -- 
    -- CP-element group 882:  join  transition  output  bypass 
    -- CP-element group 882: predecessors 
    -- CP-element group 882: 	880 
    -- CP-element group 882: 	881 
    -- CP-element group 882: successors 
    -- CP-element group 882: 	886 
    -- CP-element group 882:  members (5) 
      -- CP-element group 882: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/$exit
      -- CP-element group 882: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/$exit
      -- CP-element group 882: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/type_cast_1886/$exit
      -- CP-element group 882: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_sources/type_cast_1886/SplitProtocol/$exit
      -- CP-element group 882: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1883/phi_stmt_1883_req
      -- 
    phi_stmt_1883_req_11751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1883_req_11751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(882), ack => phi_stmt_1883_req_0); -- 
    zeropad3D_cp_element_group_882: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_882"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(880) & zeropad3D_CP_2152_elements(881);
      gj_zeropad3D_cp_element_group_882 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(882), clk => clk, reset => reset); --
    end block;
    -- CP-element group 883:  transition  input  bypass 
    -- CP-element group 883: predecessors 
    -- CP-element group 883: 	224 
    -- CP-element group 883: successors 
    -- CP-element group 883: 	885 
    -- CP-element group 883:  members (2) 
      -- CP-element group 883: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/type_cast_1882/SplitProtocol/Sample/$exit
      -- CP-element group 883: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/type_cast_1882/SplitProtocol/Sample/ra
      -- 
    ra_11768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 883_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1882_inst_ack_0, ack => zeropad3D_CP_2152_elements(883)); -- 
    -- CP-element group 884:  transition  input  bypass 
    -- CP-element group 884: predecessors 
    -- CP-element group 884: 	224 
    -- CP-element group 884: successors 
    -- CP-element group 884: 	885 
    -- CP-element group 884:  members (2) 
      -- CP-element group 884: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/type_cast_1882/SplitProtocol/Update/$exit
      -- CP-element group 884: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/type_cast_1882/SplitProtocol/Update/ca
      -- 
    ca_11773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 884_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1882_inst_ack_1, ack => zeropad3D_CP_2152_elements(884)); -- 
    -- CP-element group 885:  join  transition  output  bypass 
    -- CP-element group 885: predecessors 
    -- CP-element group 885: 	883 
    -- CP-element group 885: 	884 
    -- CP-element group 885: successors 
    -- CP-element group 885: 	886 
    -- CP-element group 885:  members (5) 
      -- CP-element group 885: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/$exit
      -- CP-element group 885: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/$exit
      -- CP-element group 885: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/type_cast_1882/$exit
      -- CP-element group 885: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_sources/type_cast_1882/SplitProtocol/$exit
      -- CP-element group 885: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/phi_stmt_1879/phi_stmt_1879_req
      -- 
    phi_stmt_1879_req_11774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1879_req_11774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(885), ack => phi_stmt_1879_req_0); -- 
    zeropad3D_cp_element_group_885: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_885"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(883) & zeropad3D_CP_2152_elements(884);
      gj_zeropad3D_cp_element_group_885 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(885), clk => clk, reset => reset); --
    end block;
    -- CP-element group 886:  join  fork  transition  place  bypass 
    -- CP-element group 886: predecessors 
    -- CP-element group 886: 	882 
    -- CP-element group 886: 	885 
    -- CP-element group 886: successors 
    -- CP-element group 886: 	887 
    -- CP-element group 886: 	888 
    -- CP-element group 886:  members (3) 
      -- CP-element group 886: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/$exit
      -- CP-element group 886: 	 branch_block_stmt_714/merge_stmt_1878_PhiReqMerge
      -- CP-element group 886: 	 branch_block_stmt_714/merge_stmt_1878_PhiAck/$entry
      -- 
    zeropad3D_cp_element_group_886: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_886"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(882) & zeropad3D_CP_2152_elements(885);
      gj_zeropad3D_cp_element_group_886 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(886), clk => clk, reset => reset); --
    end block;
    -- CP-element group 887:  transition  input  bypass 
    -- CP-element group 887: predecessors 
    -- CP-element group 887: 	886 
    -- CP-element group 887: successors 
    -- CP-element group 887: 	889 
    -- CP-element group 887:  members (1) 
      -- CP-element group 887: 	 branch_block_stmt_714/merge_stmt_1878_PhiAck/phi_stmt_1879_ack
      -- 
    phi_stmt_1879_ack_11779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 887_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1879_ack_0, ack => zeropad3D_CP_2152_elements(887)); -- 
    -- CP-element group 888:  transition  input  bypass 
    -- CP-element group 888: predecessors 
    -- CP-element group 888: 	886 
    -- CP-element group 888: successors 
    -- CP-element group 888: 	889 
    -- CP-element group 888:  members (1) 
      -- CP-element group 888: 	 branch_block_stmt_714/merge_stmt_1878_PhiAck/phi_stmt_1883_ack
      -- 
    phi_stmt_1883_ack_11780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 888_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1883_ack_0, ack => zeropad3D_CP_2152_elements(888)); -- 
    -- CP-element group 889:  join  fork  transition  place  output  bypass 
    -- CP-element group 889: predecessors 
    -- CP-element group 889: 	887 
    -- CP-element group 889: 	888 
    -- CP-element group 889: successors 
    -- CP-element group 889: 	226 
    -- CP-element group 889: 	227 
    -- CP-element group 889: 	228 
    -- CP-element group 889: 	229 
    -- CP-element group 889: 	230 
    -- CP-element group 889: 	231 
    -- CP-element group 889: 	232 
    -- CP-element group 889: 	233 
    -- CP-element group 889: 	234 
    -- CP-element group 889: 	235 
    -- CP-element group 889: 	237 
    -- CP-element group 889: 	239 
    -- CP-element group 889:  members (92) 
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011__entry__
      -- CP-element group 889: 	 branch_block_stmt_714/merge_stmt_1878__exit__
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1890_sample_start_
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1890_update_start_
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1890_Sample/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1890_Sample/rr
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1890_Update/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1890_Update/cr
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_sample_start_
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_update_start_
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_word_address_calculated
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_root_address_calculated
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Sample/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Sample/word_access_start/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Sample/word_access_start/word_0/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Sample/word_access_start/word_0/rr
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Update/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Update/word_access_complete/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Update/word_access_complete/word_0/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_pad_1899_Update/word_access_complete/word_0/cr
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_sample_start_
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_update_start_
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_word_address_calculated
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_root_address_calculated
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Sample/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Sample/word_access_start/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Sample/word_access_start/word_0/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Sample/word_access_start/word_0/rr
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Update/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Update/word_access_complete/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Update/word_access_complete/word_0/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/LOAD_depth_high_1902_Update/word_access_complete/word_0/cr
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_sample_start_
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_update_start_
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_base_address_calculated
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_word_address_calculated
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_root_address_calculated
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_base_address_resized
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_base_addr_resize/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_base_addr_resize/$exit
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_base_addr_resize/base_resize_req
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_base_addr_resize/base_resize_ack
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_base_plus_offset/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_base_plus_offset/$exit
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_base_plus_offset/sum_rename_req
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_base_plus_offset/sum_rename_ack
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_word_addrgen/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_word_addrgen/$exit
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_word_addrgen/root_register_req
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_word_addrgen/root_register_ack
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Sample/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Sample/word_access_start/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Sample/word_access_start/word_0/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Sample/word_access_start/word_0/rr
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Update/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Update/word_access_complete/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Update/word_access_complete/word_0/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1914_Update/word_access_complete/word_0/cr
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_sample_start_
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_update_start_
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_base_address_calculated
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_word_address_calculated
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_root_address_calculated
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_base_address_resized
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_base_addr_resize/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_base_addr_resize/$exit
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_base_addr_resize/base_resize_req
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_base_addr_resize/base_resize_ack
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_base_plus_offset/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_base_plus_offset/$exit
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_base_plus_offset/sum_rename_req
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_base_plus_offset/sum_rename_ack
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_word_addrgen/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_word_addrgen/$exit
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_word_addrgen/root_register_req
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_word_addrgen/root_register_ack
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Sample/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Sample/word_access_start/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Sample/word_access_start/word_0/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Sample/word_access_start/word_0/rr
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Update/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Update/word_access_complete/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Update/word_access_complete/word_0/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/ptr_deref_1926_Update/word_access_complete/word_0/cr
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1930_update_start_
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1930_Update/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1930_Update/cr
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1969_update_start_
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1969_Update/$entry
      -- CP-element group 889: 	 branch_block_stmt_714/assign_stmt_1891_to_assign_stmt_2011/type_cast_1969_Update/cr
      -- CP-element group 889: 	 branch_block_stmt_714/merge_stmt_1878_PhiAck/$exit
      -- 
    rr_4947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(889), ack => type_cast_1890_inst_req_0); -- 
    cr_4952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(889), ack => type_cast_1890_inst_req_1); -- 
    rr_4969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(889), ack => LOAD_pad_1899_load_0_req_0); -- 
    cr_4980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(889), ack => LOAD_pad_1899_load_0_req_1); -- 
    rr_5002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(889), ack => LOAD_depth_high_1902_load_0_req_0); -- 
    cr_5013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(889), ack => LOAD_depth_high_1902_load_0_req_1); -- 
    rr_5052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(889), ack => ptr_deref_1914_load_0_req_0); -- 
    cr_5063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(889), ack => ptr_deref_1914_load_0_req_1); -- 
    rr_5102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(889), ack => ptr_deref_1926_load_0_req_0); -- 
    cr_5113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(889), ack => ptr_deref_1926_load_0_req_1); -- 
    cr_5132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(889), ack => type_cast_1930_inst_req_1); -- 
    cr_5146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(889), ack => type_cast_1969_inst_req_1); -- 
    zeropad3D_cp_element_group_889: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_889"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(887) & zeropad3D_CP_2152_elements(888);
      gj_zeropad3D_cp_element_group_889 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(889), clk => clk, reset => reset); --
    end block;
    -- CP-element group 890:  transition  input  bypass 
    -- CP-element group 890: predecessors 
    -- CP-element group 890: 	3 
    -- CP-element group 890: successors 
    -- CP-element group 890: 	892 
    -- CP-element group 890:  members (2) 
      -- CP-element group 890: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/type_cast_2030/SplitProtocol/Sample/$exit
      -- CP-element group 890: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/type_cast_2030/SplitProtocol/Sample/ra
      -- 
    ra_11800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 890_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2030_inst_ack_0, ack => zeropad3D_CP_2152_elements(890)); -- 
    -- CP-element group 891:  transition  input  bypass 
    -- CP-element group 891: predecessors 
    -- CP-element group 891: 	3 
    -- CP-element group 891: successors 
    -- CP-element group 891: 	892 
    -- CP-element group 891:  members (2) 
      -- CP-element group 891: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/type_cast_2030/SplitProtocol/Update/$exit
      -- CP-element group 891: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/type_cast_2030/SplitProtocol/Update/ca
      -- 
    ca_11805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 891_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2030_inst_ack_1, ack => zeropad3D_CP_2152_elements(891)); -- 
    -- CP-element group 892:  join  transition  output  bypass 
    -- CP-element group 892: predecessors 
    -- CP-element group 892: 	890 
    -- CP-element group 892: 	891 
    -- CP-element group 892: successors 
    -- CP-element group 892: 	899 
    -- CP-element group 892:  members (5) 
      -- CP-element group 892: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/$exit
      -- CP-element group 892: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/$exit
      -- CP-element group 892: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/type_cast_2030/$exit
      -- CP-element group 892: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/type_cast_2030/SplitProtocol/$exit
      -- CP-element group 892: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_req
      -- 
    phi_stmt_2027_req_11806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2027_req_11806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(892), ack => phi_stmt_2027_req_0); -- 
    zeropad3D_cp_element_group_892: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_892"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(890) & zeropad3D_CP_2152_elements(891);
      gj_zeropad3D_cp_element_group_892 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(892), clk => clk, reset => reset); --
    end block;
    -- CP-element group 893:  transition  input  bypass 
    -- CP-element group 893: predecessors 
    -- CP-element group 893: 	3 
    -- CP-element group 893: successors 
    -- CP-element group 893: 	895 
    -- CP-element group 893:  members (2) 
      -- CP-element group 893: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Sample/$exit
      -- CP-element group 893: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Sample/ra
      -- 
    ra_11823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 893_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2017_inst_ack_0, ack => zeropad3D_CP_2152_elements(893)); -- 
    -- CP-element group 894:  transition  input  bypass 
    -- CP-element group 894: predecessors 
    -- CP-element group 894: 	3 
    -- CP-element group 894: successors 
    -- CP-element group 894: 	895 
    -- CP-element group 894:  members (2) 
      -- CP-element group 894: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Update/$exit
      -- CP-element group 894: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Update/ca
      -- 
    ca_11828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 894_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2017_inst_ack_1, ack => zeropad3D_CP_2152_elements(894)); -- 
    -- CP-element group 895:  join  transition  output  bypass 
    -- CP-element group 895: predecessors 
    -- CP-element group 895: 	893 
    -- CP-element group 895: 	894 
    -- CP-element group 895: successors 
    -- CP-element group 895: 	899 
    -- CP-element group 895:  members (5) 
      -- CP-element group 895: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/$exit
      -- CP-element group 895: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/$exit
      -- CP-element group 895: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/$exit
      -- CP-element group 895: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/$exit
      -- CP-element group 895: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_req
      -- 
    phi_stmt_2014_req_11829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2014_req_11829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(895), ack => phi_stmt_2014_req_0); -- 
    zeropad3D_cp_element_group_895: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_895"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(893) & zeropad3D_CP_2152_elements(894);
      gj_zeropad3D_cp_element_group_895 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(895), clk => clk, reset => reset); --
    end block;
    -- CP-element group 896:  transition  input  bypass 
    -- CP-element group 896: predecessors 
    -- CP-element group 896: 	3 
    -- CP-element group 896: successors 
    -- CP-element group 896: 	898 
    -- CP-element group 896:  members (2) 
      -- CP-element group 896: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2026/SplitProtocol/Sample/$exit
      -- CP-element group 896: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2026/SplitProtocol/Sample/ra
      -- 
    ra_11846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 896_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2026_inst_ack_0, ack => zeropad3D_CP_2152_elements(896)); -- 
    -- CP-element group 897:  transition  input  bypass 
    -- CP-element group 897: predecessors 
    -- CP-element group 897: 	3 
    -- CP-element group 897: successors 
    -- CP-element group 897: 	898 
    -- CP-element group 897:  members (2) 
      -- CP-element group 897: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2026/SplitProtocol/Update/$exit
      -- CP-element group 897: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2026/SplitProtocol/Update/ca
      -- 
    ca_11851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 897_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2026_inst_ack_1, ack => zeropad3D_CP_2152_elements(897)); -- 
    -- CP-element group 898:  join  transition  output  bypass 
    -- CP-element group 898: predecessors 
    -- CP-element group 898: 	896 
    -- CP-element group 898: 	897 
    -- CP-element group 898: successors 
    -- CP-element group 898: 	899 
    -- CP-element group 898:  members (5) 
      -- CP-element group 898: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/$exit
      -- CP-element group 898: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/$exit
      -- CP-element group 898: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2026/$exit
      -- CP-element group 898: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2026/SplitProtocol/$exit
      -- CP-element group 898: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_req
      -- 
    phi_stmt_2021_req_11852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2021_req_11852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(898), ack => phi_stmt_2021_req_1); -- 
    zeropad3D_cp_element_group_898: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_898"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(896) & zeropad3D_CP_2152_elements(897);
      gj_zeropad3D_cp_element_group_898 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(898), clk => clk, reset => reset); --
    end block;
    -- CP-element group 899:  join  transition  bypass 
    -- CP-element group 899: predecessors 
    -- CP-element group 899: 	892 
    -- CP-element group 899: 	895 
    -- CP-element group 899: 	898 
    -- CP-element group 899: successors 
    -- CP-element group 899: 	906 
    -- CP-element group 899:  members (1) 
      -- CP-element group 899: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_899: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_899"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(892) & zeropad3D_CP_2152_elements(895) & zeropad3D_CP_2152_elements(898);
      gj_zeropad3D_cp_element_group_899 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(899), clk => clk, reset => reset); --
    end block;
    -- CP-element group 900:  transition  output  delay-element  bypass 
    -- CP-element group 900: predecessors 
    -- CP-element group 900: 	240 
    -- CP-element group 900: successors 
    -- CP-element group 900: 	905 
    -- CP-element group 900:  members (4) 
      -- CP-element group 900: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2027/$exit
      -- CP-element group 900: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/$exit
      -- CP-element group 900: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_sources/type_cast_2033_konst_delay_trans
      -- CP-element group 900: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2027/phi_stmt_2027_req
      -- 
    phi_stmt_2027_req_11863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2027_req_11863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(900), ack => phi_stmt_2027_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(900) is a control-delay.
    cp_element_900_delay: control_delay_element  generic map(name => " 900_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(240), ack => zeropad3D_CP_2152_elements(900), clk => clk, reset =>reset);
    -- CP-element group 901:  transition  output  delay-element  bypass 
    -- CP-element group 901: predecessors 
    -- CP-element group 901: 	240 
    -- CP-element group 901: successors 
    -- CP-element group 901: 	905 
    -- CP-element group 901:  members (4) 
      -- CP-element group 901: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2014/$exit
      -- CP-element group 901: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/$exit
      -- CP-element group 901: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2020_konst_delay_trans
      -- CP-element group 901: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2014/phi_stmt_2014_req
      -- 
    phi_stmt_2014_req_11871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2014_req_11871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(901), ack => phi_stmt_2014_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(901) is a control-delay.
    cp_element_901_delay: control_delay_element  generic map(name => " 901_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(240), ack => zeropad3D_CP_2152_elements(901), clk => clk, reset =>reset);
    -- CP-element group 902:  transition  input  bypass 
    -- CP-element group 902: predecessors 
    -- CP-element group 902: 	240 
    -- CP-element group 902: successors 
    -- CP-element group 902: 	904 
    -- CP-element group 902:  members (2) 
      -- CP-element group 902: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2024/SplitProtocol/Sample/$exit
      -- CP-element group 902: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2024/SplitProtocol/Sample/ra
      -- 
    ra_11888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 902_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2024_inst_ack_0, ack => zeropad3D_CP_2152_elements(902)); -- 
    -- CP-element group 903:  transition  input  bypass 
    -- CP-element group 903: predecessors 
    -- CP-element group 903: 	240 
    -- CP-element group 903: successors 
    -- CP-element group 903: 	904 
    -- CP-element group 903:  members (2) 
      -- CP-element group 903: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2024/SplitProtocol/Update/$exit
      -- CP-element group 903: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2024/SplitProtocol/Update/ca
      -- 
    ca_11893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 903_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2024_inst_ack_1, ack => zeropad3D_CP_2152_elements(903)); -- 
    -- CP-element group 904:  join  transition  output  bypass 
    -- CP-element group 904: predecessors 
    -- CP-element group 904: 	902 
    -- CP-element group 904: 	903 
    -- CP-element group 904: successors 
    -- CP-element group 904: 	905 
    -- CP-element group 904:  members (5) 
      -- CP-element group 904: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/$exit
      -- CP-element group 904: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/$exit
      -- CP-element group 904: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2024/$exit
      -- CP-element group 904: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_sources/type_cast_2024/SplitProtocol/$exit
      -- CP-element group 904: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2021/phi_stmt_2021_req
      -- 
    phi_stmt_2021_req_11894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2021_req_11894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(904), ack => phi_stmt_2021_req_0); -- 
    zeropad3D_cp_element_group_904: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_904"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(902) & zeropad3D_CP_2152_elements(903);
      gj_zeropad3D_cp_element_group_904 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(904), clk => clk, reset => reset); --
    end block;
    -- CP-element group 905:  join  transition  bypass 
    -- CP-element group 905: predecessors 
    -- CP-element group 905: 	900 
    -- CP-element group 905: 	901 
    -- CP-element group 905: 	904 
    -- CP-element group 905: successors 
    -- CP-element group 905: 	906 
    -- CP-element group 905:  members (1) 
      -- CP-element group 905: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_905: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_905"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(900) & zeropad3D_CP_2152_elements(901) & zeropad3D_CP_2152_elements(904);
      gj_zeropad3D_cp_element_group_905 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(905), clk => clk, reset => reset); --
    end block;
    -- CP-element group 906:  merge  fork  transition  place  bypass 
    -- CP-element group 906: predecessors 
    -- CP-element group 906: 	899 
    -- CP-element group 906: 	905 
    -- CP-element group 906: successors 
    -- CP-element group 906: 	907 
    -- CP-element group 906: 	908 
    -- CP-element group 906: 	909 
    -- CP-element group 906:  members (2) 
      -- CP-element group 906: 	 branch_block_stmt_714/merge_stmt_2013_PhiReqMerge
      -- CP-element group 906: 	 branch_block_stmt_714/merge_stmt_2013_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(906) <= OrReduce(zeropad3D_CP_2152_elements(899) & zeropad3D_CP_2152_elements(905));
    -- CP-element group 907:  transition  input  bypass 
    -- CP-element group 907: predecessors 
    -- CP-element group 907: 	906 
    -- CP-element group 907: successors 
    -- CP-element group 907: 	910 
    -- CP-element group 907:  members (1) 
      -- CP-element group 907: 	 branch_block_stmt_714/merge_stmt_2013_PhiAck/phi_stmt_2014_ack
      -- 
    phi_stmt_2014_ack_11899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 907_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2014_ack_0, ack => zeropad3D_CP_2152_elements(907)); -- 
    -- CP-element group 908:  transition  input  bypass 
    -- CP-element group 908: predecessors 
    -- CP-element group 908: 	906 
    -- CP-element group 908: successors 
    -- CP-element group 908: 	910 
    -- CP-element group 908:  members (1) 
      -- CP-element group 908: 	 branch_block_stmt_714/merge_stmt_2013_PhiAck/phi_stmt_2021_ack
      -- 
    phi_stmt_2021_ack_11900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 908_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2021_ack_0, ack => zeropad3D_CP_2152_elements(908)); -- 
    -- CP-element group 909:  transition  input  bypass 
    -- CP-element group 909: predecessors 
    -- CP-element group 909: 	906 
    -- CP-element group 909: successors 
    -- CP-element group 909: 	910 
    -- CP-element group 909:  members (1) 
      -- CP-element group 909: 	 branch_block_stmt_714/merge_stmt_2013_PhiAck/phi_stmt_2027_ack
      -- 
    phi_stmt_2027_ack_11901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 909_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2027_ack_0, ack => zeropad3D_CP_2152_elements(909)); -- 
    -- CP-element group 910:  join  fork  transition  place  output  bypass 
    -- CP-element group 910: predecessors 
    -- CP-element group 910: 	907 
    -- CP-element group 910: 	908 
    -- CP-element group 910: 	909 
    -- CP-element group 910: successors 
    -- CP-element group 910: 	241 
    -- CP-element group 910: 	242 
    -- CP-element group 910:  members (10) 
      -- CP-element group 910: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046__entry__
      -- CP-element group 910: 	 branch_block_stmt_714/merge_stmt_2013__exit__
      -- CP-element group 910: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/$entry
      -- CP-element group 910: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/type_cast_2038_sample_start_
      -- CP-element group 910: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/type_cast_2038_update_start_
      -- CP-element group 910: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/type_cast_2038_Sample/$entry
      -- CP-element group 910: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/type_cast_2038_Sample/rr
      -- CP-element group 910: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/type_cast_2038_Update/$entry
      -- CP-element group 910: 	 branch_block_stmt_714/assign_stmt_2039_to_assign_stmt_2046/type_cast_2038_Update/cr
      -- CP-element group 910: 	 branch_block_stmt_714/merge_stmt_2013_PhiAck/$exit
      -- 
    rr_5158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(910), ack => type_cast_2038_inst_req_0); -- 
    cr_5163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(910), ack => type_cast_2038_inst_req_1); -- 
    zeropad3D_cp_element_group_910: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_910"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(907) & zeropad3D_CP_2152_elements(908) & zeropad3D_CP_2152_elements(909);
      gj_zeropad3D_cp_element_group_910 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(910), clk => clk, reset => reset); --
    end block;
    -- CP-element group 911:  merge  fork  transition  place  output  bypass 
    -- CP-element group 911: predecessors 
    -- CP-element group 911: 	243 
    -- CP-element group 911: 	250 
    -- CP-element group 911: 	253 
    -- CP-element group 911: 	260 
    -- CP-element group 911: successors 
    -- CP-element group 911: 	273 
    -- CP-element group 911: 	261 
    -- CP-element group 911: 	262 
    -- CP-element group 911: 	263 
    -- CP-element group 911: 	264 
    -- CP-element group 911: 	267 
    -- CP-element group 911: 	269 
    -- CP-element group 911: 	271 
    -- CP-element group 911:  members (33) 
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192__entry__
      -- CP-element group 911: 	 branch_block_stmt_714/merge_stmt_2136__exit__
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Update/word_access_complete/word_0/$entry
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Update/word_access_complete/word_0/cr
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Update/word_access_complete/$entry
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_Update/$entry
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/$entry
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2140_sample_start_
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2140_update_start_
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2140_Sample/$entry
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2140_Sample/rr
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2140_Update/$entry
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2140_Update/cr
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2145_sample_start_
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2145_update_start_
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2145_Sample/$entry
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2145_Sample/rr
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2145_Update/$entry
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2145_Update/cr
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2179_update_start_
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2179_Update/$entry
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/type_cast_2179_Update/cr
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/addr_of_2186_update_start_
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_final_index_sum_regn_update_start
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_final_index_sum_regn_Update/$entry
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/array_obj_ref_2185_final_index_sum_regn_Update/req
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/addr_of_2186_complete/$entry
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/addr_of_2186_complete/req
      -- CP-element group 911: 	 branch_block_stmt_714/assign_stmt_2141_to_assign_stmt_2192/ptr_deref_2189_update_start_
      -- CP-element group 911: 	 branch_block_stmt_714/merge_stmt_2136_PhiReqMerge
      -- CP-element group 911: 	 branch_block_stmt_714/merge_stmt_2136_PhiAck/$entry
      -- CP-element group 911: 	 branch_block_stmt_714/merge_stmt_2136_PhiAck/$exit
      -- CP-element group 911: 	 branch_block_stmt_714/merge_stmt_2136_PhiAck/dummy
      -- 
    cr_5497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(911), ack => ptr_deref_2189_store_0_req_1); -- 
    rr_5368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(911), ack => type_cast_2140_inst_req_0); -- 
    cr_5373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(911), ack => type_cast_2140_inst_req_1); -- 
    rr_5382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(911), ack => type_cast_2145_inst_req_0); -- 
    cr_5387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(911), ack => type_cast_2145_inst_req_1); -- 
    cr_5401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(911), ack => type_cast_2179_inst_req_1); -- 
    req_5432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(911), ack => array_obj_ref_2185_index_offset_req_1); -- 
    req_5447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(911), ack => addr_of_2186_final_reg_req_1); -- 
    zeropad3D_CP_2152_elements(911) <= OrReduce(zeropad3D_CP_2152_elements(243) & zeropad3D_CP_2152_elements(250) & zeropad3D_CP_2152_elements(253) & zeropad3D_CP_2152_elements(260));
    -- CP-element group 912:  merge  fork  transition  place  output  bypass 
    -- CP-element group 912: predecessors 
    -- CP-element group 912: 	274 
    -- CP-element group 912: 	294 
    -- CP-element group 912: successors 
    -- CP-element group 912: 	295 
    -- CP-element group 912: 	296 
    -- CP-element group 912:  members (13) 
      -- CP-element group 912: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319__entry__
      -- CP-element group 912: 	 branch_block_stmt_714/merge_stmt_2301__exit__
      -- CP-element group 912: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/type_cast_2305_Sample/$entry
      -- CP-element group 912: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/$entry
      -- CP-element group 912: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/type_cast_2305_sample_start_
      -- CP-element group 912: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/type_cast_2305_update_start_
      -- CP-element group 912: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/type_cast_2305_Update/cr
      -- CP-element group 912: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/type_cast_2305_Update/$entry
      -- CP-element group 912: 	 branch_block_stmt_714/assign_stmt_2306_to_assign_stmt_2319/type_cast_2305_Sample/rr
      -- CP-element group 912: 	 branch_block_stmt_714/merge_stmt_2301_PhiReqMerge
      -- CP-element group 912: 	 branch_block_stmt_714/merge_stmt_2301_PhiAck/$entry
      -- CP-element group 912: 	 branch_block_stmt_714/merge_stmt_2301_PhiAck/$exit
      -- CP-element group 912: 	 branch_block_stmt_714/merge_stmt_2301_PhiAck/dummy
      -- 
    cr_5751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(912), ack => type_cast_2305_inst_req_1); -- 
    rr_5746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(912), ack => type_cast_2305_inst_req_0); -- 
    zeropad3D_CP_2152_elements(912) <= OrReduce(zeropad3D_CP_2152_elements(274) & zeropad3D_CP_2152_elements(294));
    -- CP-element group 913:  transition  output  delay-element  bypass 
    -- CP-element group 913: predecessors 
    -- CP-element group 913: 	316 
    -- CP-element group 913: successors 
    -- CP-element group 913: 	920 
    -- CP-element group 913:  members (4) 
      -- CP-element group 913: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2420/$exit
      -- CP-element group 913: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/$exit
      -- CP-element group 913: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/type_cast_2426_konst_delay_trans
      -- CP-element group 913: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_req
      -- 
    phi_stmt_2420_req_12012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2420_req_12012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(913), ack => phi_stmt_2420_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(913) is a control-delay.
    cp_element_913_delay: control_delay_element  generic map(name => " 913_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(316), ack => zeropad3D_CP_2152_elements(913), clk => clk, reset =>reset);
    -- CP-element group 914:  transition  input  bypass 
    -- CP-element group 914: predecessors 
    -- CP-element group 914: 	316 
    -- CP-element group 914: successors 
    -- CP-element group 914: 	916 
    -- CP-element group 914:  members (2) 
      -- CP-element group 914: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2432/SplitProtocol/Sample/$exit
      -- CP-element group 914: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2432/SplitProtocol/Sample/ra
      -- 
    ra_12029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 914_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2432_inst_ack_0, ack => zeropad3D_CP_2152_elements(914)); -- 
    -- CP-element group 915:  transition  input  bypass 
    -- CP-element group 915: predecessors 
    -- CP-element group 915: 	316 
    -- CP-element group 915: successors 
    -- CP-element group 915: 	916 
    -- CP-element group 915:  members (2) 
      -- CP-element group 915: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2432/SplitProtocol/Update/$exit
      -- CP-element group 915: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2432/SplitProtocol/Update/ca
      -- 
    ca_12034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 915_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2432_inst_ack_1, ack => zeropad3D_CP_2152_elements(915)); -- 
    -- CP-element group 916:  join  transition  output  bypass 
    -- CP-element group 916: predecessors 
    -- CP-element group 916: 	914 
    -- CP-element group 916: 	915 
    -- CP-element group 916: successors 
    -- CP-element group 916: 	920 
    -- CP-element group 916:  members (5) 
      -- CP-element group 916: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/$exit
      -- CP-element group 916: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/$exit
      -- CP-element group 916: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2432/$exit
      -- CP-element group 916: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2432/SplitProtocol/$exit
      -- CP-element group 916: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_req
      -- 
    phi_stmt_2427_req_12035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2427_req_12035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(916), ack => phi_stmt_2427_req_1); -- 
    zeropad3D_cp_element_group_916: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_916"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(914) & zeropad3D_CP_2152_elements(915);
      gj_zeropad3D_cp_element_group_916 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(916), clk => clk, reset => reset); --
    end block;
    -- CP-element group 917:  transition  input  bypass 
    -- CP-element group 917: predecessors 
    -- CP-element group 917: 	316 
    -- CP-element group 917: successors 
    -- CP-element group 917: 	919 
    -- CP-element group 917:  members (2) 
      -- CP-element group 917: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Sample/$exit
      -- CP-element group 917: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Sample/ra
      -- 
    ra_12052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 917_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2438_inst_ack_0, ack => zeropad3D_CP_2152_elements(917)); -- 
    -- CP-element group 918:  transition  input  bypass 
    -- CP-element group 918: predecessors 
    -- CP-element group 918: 	316 
    -- CP-element group 918: successors 
    -- CP-element group 918: 	919 
    -- CP-element group 918:  members (2) 
      -- CP-element group 918: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Update/$exit
      -- CP-element group 918: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Update/ca
      -- 
    ca_12057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 918_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2438_inst_ack_1, ack => zeropad3D_CP_2152_elements(918)); -- 
    -- CP-element group 919:  join  transition  output  bypass 
    -- CP-element group 919: predecessors 
    -- CP-element group 919: 	917 
    -- CP-element group 919: 	918 
    -- CP-element group 919: successors 
    -- CP-element group 919: 	920 
    -- CP-element group 919:  members (5) 
      -- CP-element group 919: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/$exit
      -- CP-element group 919: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/$exit
      -- CP-element group 919: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/$exit
      -- CP-element group 919: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/$exit
      -- CP-element group 919: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_req
      -- 
    phi_stmt_2433_req_12058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2433_req_12058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(919), ack => phi_stmt_2433_req_1); -- 
    zeropad3D_cp_element_group_919: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_919"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(917) & zeropad3D_CP_2152_elements(918);
      gj_zeropad3D_cp_element_group_919 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(919), clk => clk, reset => reset); --
    end block;
    -- CP-element group 920:  join  transition  bypass 
    -- CP-element group 920: predecessors 
    -- CP-element group 920: 	913 
    -- CP-element group 920: 	916 
    -- CP-element group 920: 	919 
    -- CP-element group 920: successors 
    -- CP-element group 920: 	931 
    -- CP-element group 920:  members (1) 
      -- CP-element group 920: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_920: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_920"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(913) & zeropad3D_CP_2152_elements(916) & zeropad3D_CP_2152_elements(919);
      gj_zeropad3D_cp_element_group_920 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(920), clk => clk, reset => reset); --
    end block;
    -- CP-element group 921:  transition  input  bypass 
    -- CP-element group 921: predecessors 
    -- CP-element group 921: 	297 
    -- CP-element group 921: successors 
    -- CP-element group 921: 	923 
    -- CP-element group 921:  members (2) 
      -- CP-element group 921: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/type_cast_2423/SplitProtocol/Sample/$exit
      -- CP-element group 921: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/type_cast_2423/SplitProtocol/Sample/ra
      -- 
    ra_12078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 921_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2423_inst_ack_0, ack => zeropad3D_CP_2152_elements(921)); -- 
    -- CP-element group 922:  transition  input  bypass 
    -- CP-element group 922: predecessors 
    -- CP-element group 922: 	297 
    -- CP-element group 922: successors 
    -- CP-element group 922: 	923 
    -- CP-element group 922:  members (2) 
      -- CP-element group 922: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/type_cast_2423/SplitProtocol/Update/$exit
      -- CP-element group 922: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/type_cast_2423/SplitProtocol/Update/ca
      -- 
    ca_12083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 922_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2423_inst_ack_1, ack => zeropad3D_CP_2152_elements(922)); -- 
    -- CP-element group 923:  join  transition  output  bypass 
    -- CP-element group 923: predecessors 
    -- CP-element group 923: 	921 
    -- CP-element group 923: 	922 
    -- CP-element group 923: successors 
    -- CP-element group 923: 	930 
    -- CP-element group 923:  members (5) 
      -- CP-element group 923: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/$exit
      -- CP-element group 923: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/$exit
      -- CP-element group 923: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/type_cast_2423/$exit
      -- CP-element group 923: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_sources/type_cast_2423/SplitProtocol/$exit
      -- CP-element group 923: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2420/phi_stmt_2420_req
      -- 
    phi_stmt_2420_req_12084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2420_req_12084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(923), ack => phi_stmt_2420_req_0); -- 
    zeropad3D_cp_element_group_923: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_923"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(921) & zeropad3D_CP_2152_elements(922);
      gj_zeropad3D_cp_element_group_923 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(923), clk => clk, reset => reset); --
    end block;
    -- CP-element group 924:  transition  input  bypass 
    -- CP-element group 924: predecessors 
    -- CP-element group 924: 	297 
    -- CP-element group 924: successors 
    -- CP-element group 924: 	926 
    -- CP-element group 924:  members (2) 
      -- CP-element group 924: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2430/SplitProtocol/Sample/$exit
      -- CP-element group 924: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2430/SplitProtocol/Sample/ra
      -- 
    ra_12101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 924_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2430_inst_ack_0, ack => zeropad3D_CP_2152_elements(924)); -- 
    -- CP-element group 925:  transition  input  bypass 
    -- CP-element group 925: predecessors 
    -- CP-element group 925: 	297 
    -- CP-element group 925: successors 
    -- CP-element group 925: 	926 
    -- CP-element group 925:  members (2) 
      -- CP-element group 925: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2430/SplitProtocol/Update/$exit
      -- CP-element group 925: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2430/SplitProtocol/Update/ca
      -- 
    ca_12106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 925_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2430_inst_ack_1, ack => zeropad3D_CP_2152_elements(925)); -- 
    -- CP-element group 926:  join  transition  output  bypass 
    -- CP-element group 926: predecessors 
    -- CP-element group 926: 	924 
    -- CP-element group 926: 	925 
    -- CP-element group 926: successors 
    -- CP-element group 926: 	930 
    -- CP-element group 926:  members (5) 
      -- CP-element group 926: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/$exit
      -- CP-element group 926: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/$exit
      -- CP-element group 926: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2430/$exit
      -- CP-element group 926: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_sources/type_cast_2430/SplitProtocol/$exit
      -- CP-element group 926: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2427/phi_stmt_2427_req
      -- 
    phi_stmt_2427_req_12107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2427_req_12107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(926), ack => phi_stmt_2427_req_0); -- 
    zeropad3D_cp_element_group_926: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_926"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(924) & zeropad3D_CP_2152_elements(925);
      gj_zeropad3D_cp_element_group_926 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(926), clk => clk, reset => reset); --
    end block;
    -- CP-element group 927:  transition  input  bypass 
    -- CP-element group 927: predecessors 
    -- CP-element group 927: 	297 
    -- CP-element group 927: successors 
    -- CP-element group 927: 	929 
    -- CP-element group 927:  members (2) 
      -- CP-element group 927: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Sample/$exit
      -- CP-element group 927: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Sample/ra
      -- 
    ra_12124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 927_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2436_inst_ack_0, ack => zeropad3D_CP_2152_elements(927)); -- 
    -- CP-element group 928:  transition  input  bypass 
    -- CP-element group 928: predecessors 
    -- CP-element group 928: 	297 
    -- CP-element group 928: successors 
    -- CP-element group 928: 	929 
    -- CP-element group 928:  members (2) 
      -- CP-element group 928: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Update/$exit
      -- CP-element group 928: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Update/ca
      -- 
    ca_12129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 928_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2436_inst_ack_1, ack => zeropad3D_CP_2152_elements(928)); -- 
    -- CP-element group 929:  join  transition  output  bypass 
    -- CP-element group 929: predecessors 
    -- CP-element group 929: 	927 
    -- CP-element group 929: 	928 
    -- CP-element group 929: successors 
    -- CP-element group 929: 	930 
    -- CP-element group 929:  members (5) 
      -- CP-element group 929: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/$exit
      -- CP-element group 929: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/$exit
      -- CP-element group 929: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/$exit
      -- CP-element group 929: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/$exit
      -- CP-element group 929: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2433/phi_stmt_2433_req
      -- 
    phi_stmt_2433_req_12130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2433_req_12130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(929), ack => phi_stmt_2433_req_0); -- 
    zeropad3D_cp_element_group_929: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_929"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(927) & zeropad3D_CP_2152_elements(928);
      gj_zeropad3D_cp_element_group_929 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(929), clk => clk, reset => reset); --
    end block;
    -- CP-element group 930:  join  transition  bypass 
    -- CP-element group 930: predecessors 
    -- CP-element group 930: 	923 
    -- CP-element group 930: 	926 
    -- CP-element group 930: 	929 
    -- CP-element group 930: successors 
    -- CP-element group 930: 	931 
    -- CP-element group 930:  members (1) 
      -- CP-element group 930: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_930: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_930"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(923) & zeropad3D_CP_2152_elements(926) & zeropad3D_CP_2152_elements(929);
      gj_zeropad3D_cp_element_group_930 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(930), clk => clk, reset => reset); --
    end block;
    -- CP-element group 931:  merge  fork  transition  place  bypass 
    -- CP-element group 931: predecessors 
    -- CP-element group 931: 	920 
    -- CP-element group 931: 	930 
    -- CP-element group 931: successors 
    -- CP-element group 931: 	932 
    -- CP-element group 931: 	933 
    -- CP-element group 931: 	934 
    -- CP-element group 931:  members (2) 
      -- CP-element group 931: 	 branch_block_stmt_714/merge_stmt_2419_PhiReqMerge
      -- CP-element group 931: 	 branch_block_stmt_714/merge_stmt_2419_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(931) <= OrReduce(zeropad3D_CP_2152_elements(920) & zeropad3D_CP_2152_elements(930));
    -- CP-element group 932:  transition  input  bypass 
    -- CP-element group 932: predecessors 
    -- CP-element group 932: 	931 
    -- CP-element group 932: successors 
    -- CP-element group 932: 	935 
    -- CP-element group 932:  members (1) 
      -- CP-element group 932: 	 branch_block_stmt_714/merge_stmt_2419_PhiAck/phi_stmt_2420_ack
      -- 
    phi_stmt_2420_ack_12135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 932_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2420_ack_0, ack => zeropad3D_CP_2152_elements(932)); -- 
    -- CP-element group 933:  transition  input  bypass 
    -- CP-element group 933: predecessors 
    -- CP-element group 933: 	931 
    -- CP-element group 933: successors 
    -- CP-element group 933: 	935 
    -- CP-element group 933:  members (1) 
      -- CP-element group 933: 	 branch_block_stmt_714/merge_stmt_2419_PhiAck/phi_stmt_2427_ack
      -- 
    phi_stmt_2427_ack_12136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 933_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2427_ack_0, ack => zeropad3D_CP_2152_elements(933)); -- 
    -- CP-element group 934:  transition  input  bypass 
    -- CP-element group 934: predecessors 
    -- CP-element group 934: 	931 
    -- CP-element group 934: successors 
    -- CP-element group 934: 	935 
    -- CP-element group 934:  members (1) 
      -- CP-element group 934: 	 branch_block_stmt_714/merge_stmt_2419_PhiAck/phi_stmt_2433_ack
      -- 
    phi_stmt_2433_ack_12137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 934_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2433_ack_0, ack => zeropad3D_CP_2152_elements(934)); -- 
    -- CP-element group 935:  join  transition  bypass 
    -- CP-element group 935: predecessors 
    -- CP-element group 935: 	932 
    -- CP-element group 935: 	933 
    -- CP-element group 935: 	934 
    -- CP-element group 935: successors 
    -- CP-element group 935: 	3 
    -- CP-element group 935:  members (1) 
      -- CP-element group 935: 	 branch_block_stmt_714/merge_stmt_2419_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_935: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_935"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(932) & zeropad3D_CP_2152_elements(933) & zeropad3D_CP_2152_elements(934);
      gj_zeropad3D_cp_element_group_935 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(935), clk => clk, reset => reset); --
    end block;
    -- CP-element group 936:  transition  input  bypass 
    -- CP-element group 936: predecessors 
    -- CP-element group 936: 	315 
    -- CP-element group 936: successors 
    -- CP-element group 936: 	938 
    -- CP-element group 936:  members (2) 
      -- CP-element group 936: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/type_cast_2445/SplitProtocol/Sample/$exit
      -- CP-element group 936: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/type_cast_2445/SplitProtocol/Sample/ra
      -- 
    ra_12157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 936_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2445_inst_ack_0, ack => zeropad3D_CP_2152_elements(936)); -- 
    -- CP-element group 937:  transition  input  bypass 
    -- CP-element group 937: predecessors 
    -- CP-element group 937: 	315 
    -- CP-element group 937: successors 
    -- CP-element group 937: 	938 
    -- CP-element group 937:  members (2) 
      -- CP-element group 937: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/type_cast_2445/SplitProtocol/Update/$exit
      -- CP-element group 937: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/type_cast_2445/SplitProtocol/Update/ca
      -- 
    ca_12162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 937_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2445_inst_ack_1, ack => zeropad3D_CP_2152_elements(937)); -- 
    -- CP-element group 938:  join  transition  output  bypass 
    -- CP-element group 938: predecessors 
    -- CP-element group 938: 	936 
    -- CP-element group 938: 	937 
    -- CP-element group 938: successors 
    -- CP-element group 938: 	945 
    -- CP-element group 938:  members (5) 
      -- CP-element group 938: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/$exit
      -- CP-element group 938: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/$exit
      -- CP-element group 938: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/type_cast_2445/$exit
      -- CP-element group 938: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_sources/type_cast_2445/SplitProtocol/$exit
      -- CP-element group 938: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2442/phi_stmt_2442_req
      -- 
    phi_stmt_2442_req_12163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2442_req_12163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(938), ack => phi_stmt_2442_req_0); -- 
    zeropad3D_cp_element_group_938: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_938"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(936) & zeropad3D_CP_2152_elements(937);
      gj_zeropad3D_cp_element_group_938 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(938), clk => clk, reset => reset); --
    end block;
    -- CP-element group 939:  transition  input  bypass 
    -- CP-element group 939: predecessors 
    -- CP-element group 939: 	315 
    -- CP-element group 939: successors 
    -- CP-element group 939: 	941 
    -- CP-element group 939:  members (2) 
      -- CP-element group 939: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Sample/$exit
      -- CP-element group 939: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Sample/ra
      -- 
    ra_12180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 939_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2449_inst_ack_0, ack => zeropad3D_CP_2152_elements(939)); -- 
    -- CP-element group 940:  transition  input  bypass 
    -- CP-element group 940: predecessors 
    -- CP-element group 940: 	315 
    -- CP-element group 940: successors 
    -- CP-element group 940: 	941 
    -- CP-element group 940:  members (2) 
      -- CP-element group 940: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Update/$exit
      -- CP-element group 940: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Update/ca
      -- 
    ca_12185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 940_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2449_inst_ack_1, ack => zeropad3D_CP_2152_elements(940)); -- 
    -- CP-element group 941:  join  transition  output  bypass 
    -- CP-element group 941: predecessors 
    -- CP-element group 941: 	939 
    -- CP-element group 941: 	940 
    -- CP-element group 941: successors 
    -- CP-element group 941: 	945 
    -- CP-element group 941:  members (5) 
      -- CP-element group 941: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/$exit
      -- CP-element group 941: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/$exit
      -- CP-element group 941: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/$exit
      -- CP-element group 941: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/$exit
      -- CP-element group 941: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2446/phi_stmt_2446_req
      -- 
    phi_stmt_2446_req_12186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2446_req_12186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(941), ack => phi_stmt_2446_req_0); -- 
    zeropad3D_cp_element_group_941: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_941"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(939) & zeropad3D_CP_2152_elements(940);
      gj_zeropad3D_cp_element_group_941 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(941), clk => clk, reset => reset); --
    end block;
    -- CP-element group 942:  transition  input  bypass 
    -- CP-element group 942: predecessors 
    -- CP-element group 942: 	315 
    -- CP-element group 942: successors 
    -- CP-element group 942: 	944 
    -- CP-element group 942:  members (2) 
      -- CP-element group 942: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/type_cast_2453/SplitProtocol/Sample/$exit
      -- CP-element group 942: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/type_cast_2453/SplitProtocol/Sample/ra
      -- 
    ra_12203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 942_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2453_inst_ack_0, ack => zeropad3D_CP_2152_elements(942)); -- 
    -- CP-element group 943:  transition  input  bypass 
    -- CP-element group 943: predecessors 
    -- CP-element group 943: 	315 
    -- CP-element group 943: successors 
    -- CP-element group 943: 	944 
    -- CP-element group 943:  members (2) 
      -- CP-element group 943: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/type_cast_2453/SplitProtocol/Update/$exit
      -- CP-element group 943: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/type_cast_2453/SplitProtocol/Update/ca
      -- 
    ca_12208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 943_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2453_inst_ack_1, ack => zeropad3D_CP_2152_elements(943)); -- 
    -- CP-element group 944:  join  transition  output  bypass 
    -- CP-element group 944: predecessors 
    -- CP-element group 944: 	942 
    -- CP-element group 944: 	943 
    -- CP-element group 944: successors 
    -- CP-element group 944: 	945 
    -- CP-element group 944:  members (5) 
      -- CP-element group 944: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/$exit
      -- CP-element group 944: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/$exit
      -- CP-element group 944: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/type_cast_2453/$exit
      -- CP-element group 944: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_sources/type_cast_2453/SplitProtocol/$exit
      -- CP-element group 944: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/phi_stmt_2450/phi_stmt_2450_req
      -- 
    phi_stmt_2450_req_12209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2450_req_12209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(944), ack => phi_stmt_2450_req_0); -- 
    zeropad3D_cp_element_group_944: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_944"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(942) & zeropad3D_CP_2152_elements(943);
      gj_zeropad3D_cp_element_group_944 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(944), clk => clk, reset => reset); --
    end block;
    -- CP-element group 945:  join  fork  transition  place  bypass 
    -- CP-element group 945: predecessors 
    -- CP-element group 945: 	938 
    -- CP-element group 945: 	941 
    -- CP-element group 945: 	944 
    -- CP-element group 945: successors 
    -- CP-element group 945: 	946 
    -- CP-element group 945: 	947 
    -- CP-element group 945: 	948 
    -- CP-element group 945:  members (3) 
      -- CP-element group 945: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/$exit
      -- CP-element group 945: 	 branch_block_stmt_714/merge_stmt_2441_PhiReqMerge
      -- CP-element group 945: 	 branch_block_stmt_714/merge_stmt_2441_PhiAck/$entry
      -- 
    zeropad3D_cp_element_group_945: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_945"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(938) & zeropad3D_CP_2152_elements(941) & zeropad3D_CP_2152_elements(944);
      gj_zeropad3D_cp_element_group_945 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(945), clk => clk, reset => reset); --
    end block;
    -- CP-element group 946:  transition  input  bypass 
    -- CP-element group 946: predecessors 
    -- CP-element group 946: 	945 
    -- CP-element group 946: successors 
    -- CP-element group 946: 	949 
    -- CP-element group 946:  members (1) 
      -- CP-element group 946: 	 branch_block_stmt_714/merge_stmt_2441_PhiAck/phi_stmt_2442_ack
      -- 
    phi_stmt_2442_ack_12214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 946_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2442_ack_0, ack => zeropad3D_CP_2152_elements(946)); -- 
    -- CP-element group 947:  transition  input  bypass 
    -- CP-element group 947: predecessors 
    -- CP-element group 947: 	945 
    -- CP-element group 947: successors 
    -- CP-element group 947: 	949 
    -- CP-element group 947:  members (1) 
      -- CP-element group 947: 	 branch_block_stmt_714/merge_stmt_2441_PhiAck/phi_stmt_2446_ack
      -- 
    phi_stmt_2446_ack_12215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 947_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2446_ack_0, ack => zeropad3D_CP_2152_elements(947)); -- 
    -- CP-element group 948:  transition  input  bypass 
    -- CP-element group 948: predecessors 
    -- CP-element group 948: 	945 
    -- CP-element group 948: successors 
    -- CP-element group 948: 	949 
    -- CP-element group 948:  members (1) 
      -- CP-element group 948: 	 branch_block_stmt_714/merge_stmt_2441_PhiAck/phi_stmt_2450_ack
      -- 
    phi_stmt_2450_ack_12216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 948_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2450_ack_0, ack => zeropad3D_CP_2152_elements(948)); -- 
    -- CP-element group 949:  join  fork  transition  place  output  bypass 
    -- CP-element group 949: predecessors 
    -- CP-element group 949: 	946 
    -- CP-element group 949: 	947 
    -- CP-element group 949: 	948 
    -- CP-element group 949: successors 
    -- CP-element group 949: 	317 
    -- CP-element group 949: 	318 
    -- CP-element group 949: 	319 
    -- CP-element group 949: 	320 
    -- CP-element group 949: 	321 
    -- CP-element group 949: 	322 
    -- CP-element group 949: 	323 
    -- CP-element group 949: 	324 
    -- CP-element group 949: 	325 
    -- CP-element group 949: 	327 
    -- CP-element group 949: 	326 
    -- CP-element group 949: 	328 
    -- CP-element group 949: 	330 
    -- CP-element group 949: 	332 
    -- CP-element group 949:  members (98) 
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588__entry__
      -- CP-element group 949: 	 branch_block_stmt_714/merge_stmt_2441__exit__
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2457_sample_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2457_update_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2457_Sample/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2457_Sample/rr
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2457_Update/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2457_Update/cr
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2467_sample_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2467_update_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2467_Sample/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2467_Sample/rr
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2467_Update/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2467_Update/cr
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_sample_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_update_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_word_address_calculated
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_root_address_calculated
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Sample/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Sample/word_access_start/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Sample/word_access_start/word_0/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Sample/word_access_start/word_0/rr
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Update/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Update/word_access_complete/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Update/word_access_complete/word_0/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_pad_2476_Update/word_access_complete/word_0/cr
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_sample_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_update_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_word_address_calculated
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_root_address_calculated
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Sample/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Sample/word_access_start/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Sample/word_access_start/word_0/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Sample/word_access_start/word_0/rr
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Update/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Update/word_access_complete/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Update/word_access_complete/word_0/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/LOAD_depth_high_2479_Update/word_access_complete/word_0/cr
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_sample_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_update_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_base_address_calculated
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_word_address_calculated
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_root_address_calculated
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_base_address_resized
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_base_addr_resize/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_base_addr_resize/$exit
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_base_addr_resize/base_resize_req
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_base_addr_resize/base_resize_ack
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_base_plus_offset/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_base_plus_offset/$exit
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_base_plus_offset/sum_rename_req
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_base_plus_offset/sum_rename_ack
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_word_addrgen/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_word_addrgen/$exit
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_word_addrgen/root_register_req
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_word_addrgen/root_register_ack
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Sample/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Sample/word_access_start/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Sample/word_access_start/word_0/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Sample/word_access_start/word_0/rr
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Update/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Update/word_access_complete/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Update/word_access_complete/word_0/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2491_Update/word_access_complete/word_0/cr
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_sample_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_update_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_base_address_calculated
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_word_address_calculated
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_root_address_calculated
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_base_address_resized
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_base_addr_resize/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_base_addr_resize/$exit
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_base_addr_resize/base_resize_req
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_base_addr_resize/base_resize_ack
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_base_plus_offset/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_base_plus_offset/$exit
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_base_plus_offset/sum_rename_req
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_base_plus_offset/sum_rename_ack
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_word_addrgen/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_word_addrgen/$exit
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_word_addrgen/root_register_req
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_word_addrgen/root_register_ack
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Sample/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Sample/word_access_start/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Sample/word_access_start/word_0/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Sample/word_access_start/word_0/rr
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Update/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Update/word_access_complete/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Update/word_access_complete/word_0/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/ptr_deref_2503_Update/word_access_complete/word_0/cr
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2507_update_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2507_Update/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2507_Update/cr
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2546_update_start_
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2546_Update/$entry
      -- CP-element group 949: 	 branch_block_stmt_714/assign_stmt_2458_to_assign_stmt_2588/type_cast_2546_Update/cr
      -- CP-element group 949: 	 branch_block_stmt_714/merge_stmt_2441_PhiAck/$exit
      -- 
    rr_5943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => type_cast_2457_inst_req_0); -- 
    cr_5948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => type_cast_2457_inst_req_1); -- 
    rr_5957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => type_cast_2467_inst_req_0); -- 
    cr_5962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => type_cast_2467_inst_req_1); -- 
    rr_5979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => LOAD_pad_2476_load_0_req_0); -- 
    cr_5990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => LOAD_pad_2476_load_0_req_1); -- 
    rr_6012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => LOAD_depth_high_2479_load_0_req_0); -- 
    cr_6023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => LOAD_depth_high_2479_load_0_req_1); -- 
    rr_6062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => ptr_deref_2491_load_0_req_0); -- 
    cr_6073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => ptr_deref_2491_load_0_req_1); -- 
    rr_6112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => ptr_deref_2503_load_0_req_0); -- 
    cr_6123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => ptr_deref_2503_load_0_req_1); -- 
    cr_6142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => type_cast_2507_inst_req_1); -- 
    cr_6156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => type_cast_2546_inst_req_1); -- 
    zeropad3D_cp_element_group_949: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_949"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(946) & zeropad3D_CP_2152_elements(947) & zeropad3D_CP_2152_elements(948);
      gj_zeropad3D_cp_element_group_949 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(949), clk => clk, reset => reset); --
    end block;
    -- CP-element group 950:  transition  input  bypass 
    -- CP-element group 950: predecessors 
    -- CP-element group 950: 	4 
    -- CP-element group 950: successors 
    -- CP-element group 950: 	952 
    -- CP-element group 950:  members (2) 
      -- CP-element group 950: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/type_cast_2597/SplitProtocol/Sample/$exit
      -- CP-element group 950: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/type_cast_2597/SplitProtocol/Sample/ra
      -- 
    ra_12236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 950_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2597_inst_ack_0, ack => zeropad3D_CP_2152_elements(950)); -- 
    -- CP-element group 951:  transition  input  bypass 
    -- CP-element group 951: predecessors 
    -- CP-element group 951: 	4 
    -- CP-element group 951: successors 
    -- CP-element group 951: 	952 
    -- CP-element group 951:  members (2) 
      -- CP-element group 951: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/type_cast_2597/SplitProtocol/Update/$exit
      -- CP-element group 951: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/type_cast_2597/SplitProtocol/Update/ca
      -- 
    ca_12241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 951_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2597_inst_ack_1, ack => zeropad3D_CP_2152_elements(951)); -- 
    -- CP-element group 952:  join  transition  output  bypass 
    -- CP-element group 952: predecessors 
    -- CP-element group 952: 	950 
    -- CP-element group 952: 	951 
    -- CP-element group 952: successors 
    -- CP-element group 952: 	959 
    -- CP-element group 952:  members (5) 
      -- CP-element group 952: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/$exit
      -- CP-element group 952: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/$exit
      -- CP-element group 952: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/type_cast_2597/$exit
      -- CP-element group 952: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/type_cast_2597/SplitProtocol/$exit
      -- CP-element group 952: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_req
      -- 
    phi_stmt_2591_req_12242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2591_req_12242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(952), ack => phi_stmt_2591_req_1); -- 
    zeropad3D_cp_element_group_952: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_952"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(950) & zeropad3D_CP_2152_elements(951);
      gj_zeropad3D_cp_element_group_952 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(952), clk => clk, reset => reset); --
    end block;
    -- CP-element group 953:  transition  input  bypass 
    -- CP-element group 953: predecessors 
    -- CP-element group 953: 	4 
    -- CP-element group 953: successors 
    -- CP-element group 953: 	955 
    -- CP-element group 953:  members (2) 
      -- CP-element group 953: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2603/SplitProtocol/Sample/$exit
      -- CP-element group 953: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2603/SplitProtocol/Sample/ra
      -- 
    ra_12259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 953_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2603_inst_ack_0, ack => zeropad3D_CP_2152_elements(953)); -- 
    -- CP-element group 954:  transition  input  bypass 
    -- CP-element group 954: predecessors 
    -- CP-element group 954: 	4 
    -- CP-element group 954: successors 
    -- CP-element group 954: 	955 
    -- CP-element group 954:  members (2) 
      -- CP-element group 954: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2603/SplitProtocol/Update/$exit
      -- CP-element group 954: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2603/SplitProtocol/Update/ca
      -- 
    ca_12264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 954_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2603_inst_ack_1, ack => zeropad3D_CP_2152_elements(954)); -- 
    -- CP-element group 955:  join  transition  output  bypass 
    -- CP-element group 955: predecessors 
    -- CP-element group 955: 	953 
    -- CP-element group 955: 	954 
    -- CP-element group 955: successors 
    -- CP-element group 955: 	959 
    -- CP-element group 955:  members (5) 
      -- CP-element group 955: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/$exit
      -- CP-element group 955: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/$exit
      -- CP-element group 955: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2603/$exit
      -- CP-element group 955: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2603/SplitProtocol/$exit
      -- CP-element group 955: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_req
      -- 
    phi_stmt_2598_req_12265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2598_req_12265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(955), ack => phi_stmt_2598_req_1); -- 
    zeropad3D_cp_element_group_955: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_955"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(953) & zeropad3D_CP_2152_elements(954);
      gj_zeropad3D_cp_element_group_955 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(955), clk => clk, reset => reset); --
    end block;
    -- CP-element group 956:  transition  input  bypass 
    -- CP-element group 956: predecessors 
    -- CP-element group 956: 	4 
    -- CP-element group 956: successors 
    -- CP-element group 956: 	958 
    -- CP-element group 956:  members (2) 
      -- CP-element group 956: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2609/SplitProtocol/Sample/$exit
      -- CP-element group 956: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2609/SplitProtocol/Sample/ra
      -- 
    ra_12282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 956_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2609_inst_ack_0, ack => zeropad3D_CP_2152_elements(956)); -- 
    -- CP-element group 957:  transition  input  bypass 
    -- CP-element group 957: predecessors 
    -- CP-element group 957: 	4 
    -- CP-element group 957: successors 
    -- CP-element group 957: 	958 
    -- CP-element group 957:  members (2) 
      -- CP-element group 957: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2609/SplitProtocol/Update/$exit
      -- CP-element group 957: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2609/SplitProtocol/Update/ca
      -- 
    ca_12287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 957_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2609_inst_ack_1, ack => zeropad3D_CP_2152_elements(957)); -- 
    -- CP-element group 958:  join  transition  output  bypass 
    -- CP-element group 958: predecessors 
    -- CP-element group 958: 	956 
    -- CP-element group 958: 	957 
    -- CP-element group 958: successors 
    -- CP-element group 958: 	959 
    -- CP-element group 958:  members (5) 
      -- CP-element group 958: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/$exit
      -- CP-element group 958: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/$exit
      -- CP-element group 958: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2609/$exit
      -- CP-element group 958: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2609/SplitProtocol/$exit
      -- CP-element group 958: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_req
      -- 
    phi_stmt_2604_req_12288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2604_req_12288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(958), ack => phi_stmt_2604_req_1); -- 
    zeropad3D_cp_element_group_958: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_958"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(956) & zeropad3D_CP_2152_elements(957);
      gj_zeropad3D_cp_element_group_958 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(958), clk => clk, reset => reset); --
    end block;
    -- CP-element group 959:  join  transition  bypass 
    -- CP-element group 959: predecessors 
    -- CP-element group 959: 	952 
    -- CP-element group 959: 	955 
    -- CP-element group 959: 	958 
    -- CP-element group 959: successors 
    -- CP-element group 959: 	968 
    -- CP-element group 959:  members (1) 
      -- CP-element group 959: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_959: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_959"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(952) & zeropad3D_CP_2152_elements(955) & zeropad3D_CP_2152_elements(958);
      gj_zeropad3D_cp_element_group_959 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(959), clk => clk, reset => reset); --
    end block;
    -- CP-element group 960:  transition  output  delay-element  bypass 
    -- CP-element group 960: predecessors 
    -- CP-element group 960: 	333 
    -- CP-element group 960: successors 
    -- CP-element group 960: 	967 
    -- CP-element group 960:  members (4) 
      -- CP-element group 960: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2591/$exit
      -- CP-element group 960: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/$exit
      -- CP-element group 960: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_sources/type_cast_2595_konst_delay_trans
      -- CP-element group 960: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2591/phi_stmt_2591_req
      -- 
    phi_stmt_2591_req_12299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2591_req_12299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(960), ack => phi_stmt_2591_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(960) is a control-delay.
    cp_element_960_delay: control_delay_element  generic map(name => " 960_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(333), ack => zeropad3D_CP_2152_elements(960), clk => clk, reset =>reset);
    -- CP-element group 961:  transition  input  bypass 
    -- CP-element group 961: predecessors 
    -- CP-element group 961: 	333 
    -- CP-element group 961: successors 
    -- CP-element group 961: 	963 
    -- CP-element group 961:  members (2) 
      -- CP-element group 961: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2601/SplitProtocol/Sample/$exit
      -- CP-element group 961: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2601/SplitProtocol/Sample/ra
      -- 
    ra_12316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 961_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2601_inst_ack_0, ack => zeropad3D_CP_2152_elements(961)); -- 
    -- CP-element group 962:  transition  input  bypass 
    -- CP-element group 962: predecessors 
    -- CP-element group 962: 	333 
    -- CP-element group 962: successors 
    -- CP-element group 962: 	963 
    -- CP-element group 962:  members (2) 
      -- CP-element group 962: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2601/SplitProtocol/Update/$exit
      -- CP-element group 962: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2601/SplitProtocol/Update/ca
      -- 
    ca_12321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 962_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2601_inst_ack_1, ack => zeropad3D_CP_2152_elements(962)); -- 
    -- CP-element group 963:  join  transition  output  bypass 
    -- CP-element group 963: predecessors 
    -- CP-element group 963: 	961 
    -- CP-element group 963: 	962 
    -- CP-element group 963: successors 
    -- CP-element group 963: 	967 
    -- CP-element group 963:  members (5) 
      -- CP-element group 963: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/$exit
      -- CP-element group 963: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/$exit
      -- CP-element group 963: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2601/$exit
      -- CP-element group 963: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_sources/type_cast_2601/SplitProtocol/$exit
      -- CP-element group 963: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2598/phi_stmt_2598_req
      -- 
    phi_stmt_2598_req_12322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2598_req_12322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(963), ack => phi_stmt_2598_req_0); -- 
    zeropad3D_cp_element_group_963: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_963"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(961) & zeropad3D_CP_2152_elements(962);
      gj_zeropad3D_cp_element_group_963 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(963), clk => clk, reset => reset); --
    end block;
    -- CP-element group 964:  transition  input  bypass 
    -- CP-element group 964: predecessors 
    -- CP-element group 964: 	333 
    -- CP-element group 964: successors 
    -- CP-element group 964: 	966 
    -- CP-element group 964:  members (2) 
      -- CP-element group 964: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Sample/$exit
      -- CP-element group 964: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Sample/ra
      -- 
    ra_12339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 964_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2607_inst_ack_0, ack => zeropad3D_CP_2152_elements(964)); -- 
    -- CP-element group 965:  transition  input  bypass 
    -- CP-element group 965: predecessors 
    -- CP-element group 965: 	333 
    -- CP-element group 965: successors 
    -- CP-element group 965: 	966 
    -- CP-element group 965:  members (2) 
      -- CP-element group 965: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Update/$exit
      -- CP-element group 965: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Update/ca
      -- 
    ca_12344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 965_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2607_inst_ack_1, ack => zeropad3D_CP_2152_elements(965)); -- 
    -- CP-element group 966:  join  transition  output  bypass 
    -- CP-element group 966: predecessors 
    -- CP-element group 966: 	964 
    -- CP-element group 966: 	965 
    -- CP-element group 966: successors 
    -- CP-element group 966: 	967 
    -- CP-element group 966:  members (5) 
      -- CP-element group 966: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/$exit
      -- CP-element group 966: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/$exit
      -- CP-element group 966: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/$exit
      -- CP-element group 966: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/$exit
      -- CP-element group 966: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2604/phi_stmt_2604_req
      -- 
    phi_stmt_2604_req_12345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2604_req_12345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(966), ack => phi_stmt_2604_req_0); -- 
    zeropad3D_cp_element_group_966: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_966"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(964) & zeropad3D_CP_2152_elements(965);
      gj_zeropad3D_cp_element_group_966 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(966), clk => clk, reset => reset); --
    end block;
    -- CP-element group 967:  join  transition  bypass 
    -- CP-element group 967: predecessors 
    -- CP-element group 967: 	960 
    -- CP-element group 967: 	963 
    -- CP-element group 967: 	966 
    -- CP-element group 967: successors 
    -- CP-element group 967: 	968 
    -- CP-element group 967:  members (1) 
      -- CP-element group 967: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_967: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_967"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(960) & zeropad3D_CP_2152_elements(963) & zeropad3D_CP_2152_elements(966);
      gj_zeropad3D_cp_element_group_967 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(967), clk => clk, reset => reset); --
    end block;
    -- CP-element group 968:  merge  fork  transition  place  bypass 
    -- CP-element group 968: predecessors 
    -- CP-element group 968: 	959 
    -- CP-element group 968: 	967 
    -- CP-element group 968: successors 
    -- CP-element group 968: 	969 
    -- CP-element group 968: 	970 
    -- CP-element group 968: 	971 
    -- CP-element group 968:  members (2) 
      -- CP-element group 968: 	 branch_block_stmt_714/merge_stmt_2590_PhiReqMerge
      -- CP-element group 968: 	 branch_block_stmt_714/merge_stmt_2590_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(968) <= OrReduce(zeropad3D_CP_2152_elements(959) & zeropad3D_CP_2152_elements(967));
    -- CP-element group 969:  transition  input  bypass 
    -- CP-element group 969: predecessors 
    -- CP-element group 969: 	968 
    -- CP-element group 969: successors 
    -- CP-element group 969: 	972 
    -- CP-element group 969:  members (1) 
      -- CP-element group 969: 	 branch_block_stmt_714/merge_stmt_2590_PhiAck/phi_stmt_2591_ack
      -- 
    phi_stmt_2591_ack_12350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 969_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2591_ack_0, ack => zeropad3D_CP_2152_elements(969)); -- 
    -- CP-element group 970:  transition  input  bypass 
    -- CP-element group 970: predecessors 
    -- CP-element group 970: 	968 
    -- CP-element group 970: successors 
    -- CP-element group 970: 	972 
    -- CP-element group 970:  members (1) 
      -- CP-element group 970: 	 branch_block_stmt_714/merge_stmt_2590_PhiAck/phi_stmt_2598_ack
      -- 
    phi_stmt_2598_ack_12351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 970_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2598_ack_0, ack => zeropad3D_CP_2152_elements(970)); -- 
    -- CP-element group 971:  transition  input  bypass 
    -- CP-element group 971: predecessors 
    -- CP-element group 971: 	968 
    -- CP-element group 971: successors 
    -- CP-element group 971: 	972 
    -- CP-element group 971:  members (1) 
      -- CP-element group 971: 	 branch_block_stmt_714/merge_stmt_2590_PhiAck/phi_stmt_2604_ack
      -- 
    phi_stmt_2604_ack_12352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 971_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2604_ack_0, ack => zeropad3D_CP_2152_elements(971)); -- 
    -- CP-element group 972:  join  fork  transition  place  output  bypass 
    -- CP-element group 972: predecessors 
    -- CP-element group 972: 	969 
    -- CP-element group 972: 	970 
    -- CP-element group 972: 	971 
    -- CP-element group 972: successors 
    -- CP-element group 972: 	334 
    -- CP-element group 972: 	335 
    -- CP-element group 972:  members (10) 
      -- CP-element group 972: 	 branch_block_stmt_714/merge_stmt_2590__exit__
      -- CP-element group 972: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622__entry__
      -- CP-element group 972: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/$entry
      -- CP-element group 972: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/type_cast_2614_sample_start_
      -- CP-element group 972: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/type_cast_2614_update_start_
      -- CP-element group 972: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/type_cast_2614_Sample/$entry
      -- CP-element group 972: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/type_cast_2614_Sample/rr
      -- CP-element group 972: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/type_cast_2614_Update/$entry
      -- CP-element group 972: 	 branch_block_stmt_714/assign_stmt_2615_to_assign_stmt_2622/type_cast_2614_Update/cr
      -- CP-element group 972: 	 branch_block_stmt_714/merge_stmt_2590_PhiAck/$exit
      -- 
    rr_6168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(972), ack => type_cast_2614_inst_req_0); -- 
    cr_6173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(972), ack => type_cast_2614_inst_req_1); -- 
    zeropad3D_cp_element_group_972: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_972"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(969) & zeropad3D_CP_2152_elements(970) & zeropad3D_CP_2152_elements(971);
      gj_zeropad3D_cp_element_group_972 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(972), clk => clk, reset => reset); --
    end block;
    -- CP-element group 973:  merge  fork  transition  place  output  bypass 
    -- CP-element group 973: predecessors 
    -- CP-element group 973: 	336 
    -- CP-element group 973: 	343 
    -- CP-element group 973: 	346 
    -- CP-element group 973: 	353 
    -- CP-element group 973: successors 
    -- CP-element group 973: 	354 
    -- CP-element group 973: 	355 
    -- CP-element group 973: 	356 
    -- CP-element group 973: 	357 
    -- CP-element group 973: 	360 
    -- CP-element group 973: 	362 
    -- CP-element group 973: 	364 
    -- CP-element group 973: 	366 
    -- CP-element group 973:  members (33) 
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762__entry__
      -- CP-element group 973: 	 branch_block_stmt_714/merge_stmt_2706__exit__
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/$entry
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2710_sample_start_
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2710_update_start_
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2710_Sample/$entry
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2710_Sample/rr
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2710_Update/$entry
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2710_Update/cr
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2715_sample_start_
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2715_update_start_
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2715_Sample/$entry
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2715_Sample/rr
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2715_Update/$entry
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2715_Update/cr
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2749_update_start_
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2749_Update/$entry
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/type_cast_2749_Update/cr
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/addr_of_2756_update_start_
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_final_index_sum_regn_update_start
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_final_index_sum_regn_Update/$entry
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/array_obj_ref_2755_final_index_sum_regn_Update/req
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/addr_of_2756_complete/$entry
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/addr_of_2756_complete/req
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_update_start_
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Update/$entry
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Update/word_access_complete/$entry
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Update/word_access_complete/word_0/$entry
      -- CP-element group 973: 	 branch_block_stmt_714/assign_stmt_2711_to_assign_stmt_2762/ptr_deref_2759_Update/word_access_complete/word_0/cr
      -- CP-element group 973: 	 branch_block_stmt_714/merge_stmt_2706_PhiReqMerge
      -- CP-element group 973: 	 branch_block_stmt_714/merge_stmt_2706_PhiAck/$entry
      -- CP-element group 973: 	 branch_block_stmt_714/merge_stmt_2706_PhiAck/$exit
      -- CP-element group 973: 	 branch_block_stmt_714/merge_stmt_2706_PhiAck/dummy
      -- 
    rr_6378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(973), ack => type_cast_2710_inst_req_0); -- 
    cr_6383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(973), ack => type_cast_2710_inst_req_1); -- 
    rr_6392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(973), ack => type_cast_2715_inst_req_0); -- 
    cr_6397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(973), ack => type_cast_2715_inst_req_1); -- 
    cr_6411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(973), ack => type_cast_2749_inst_req_1); -- 
    req_6442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(973), ack => array_obj_ref_2755_index_offset_req_1); -- 
    req_6457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(973), ack => addr_of_2756_final_reg_req_1); -- 
    cr_6507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(973), ack => ptr_deref_2759_store_0_req_1); -- 
    zeropad3D_CP_2152_elements(973) <= OrReduce(zeropad3D_CP_2152_elements(336) & zeropad3D_CP_2152_elements(343) & zeropad3D_CP_2152_elements(346) & zeropad3D_CP_2152_elements(353));
    -- CP-element group 974:  merge  fork  transition  place  output  bypass 
    -- CP-element group 974: predecessors 
    -- CP-element group 974: 	367 
    -- CP-element group 974: 	387 
    -- CP-element group 974: successors 
    -- CP-element group 974: 	388 
    -- CP-element group 974: 	389 
    -- CP-element group 974:  members (13) 
      -- CP-element group 974: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889__entry__
      -- CP-element group 974: 	 branch_block_stmt_714/merge_stmt_2871__exit__
      -- CP-element group 974: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/type_cast_2875_Update/cr
      -- CP-element group 974: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/type_cast_2875_Update/$entry
      -- CP-element group 974: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/type_cast_2875_Sample/rr
      -- CP-element group 974: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/type_cast_2875_Sample/$entry
      -- CP-element group 974: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/type_cast_2875_update_start_
      -- CP-element group 974: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/type_cast_2875_sample_start_
      -- CP-element group 974: 	 branch_block_stmt_714/assign_stmt_2876_to_assign_stmt_2889/$entry
      -- CP-element group 974: 	 branch_block_stmt_714/merge_stmt_2871_PhiReqMerge
      -- CP-element group 974: 	 branch_block_stmt_714/merge_stmt_2871_PhiAck/$entry
      -- CP-element group 974: 	 branch_block_stmt_714/merge_stmt_2871_PhiAck/$exit
      -- CP-element group 974: 	 branch_block_stmt_714/merge_stmt_2871_PhiAck/dummy
      -- 
    cr_6761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(974), ack => type_cast_2875_inst_req_1); -- 
    rr_6756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(974), ack => type_cast_2875_inst_req_0); -- 
    zeropad3D_CP_2152_elements(974) <= OrReduce(zeropad3D_CP_2152_elements(367) & zeropad3D_CP_2152_elements(387));
    -- CP-element group 975:  transition  output  delay-element  bypass 
    -- CP-element group 975: predecessors 
    -- CP-element group 975: 	409 
    -- CP-element group 975: successors 
    -- CP-element group 975: 	982 
    -- CP-element group 975:  members (4) 
      -- CP-element group 975: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_req
      -- CP-element group 975: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/type_cast_2989_konst_delay_trans
      -- CP-element group 975: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/$exit
      -- CP-element group 975: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2983/$exit
      -- 
    phi_stmt_2983_req_12463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2983_req_12463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(975), ack => phi_stmt_2983_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(975) is a control-delay.
    cp_element_975_delay: control_delay_element  generic map(name => " 975_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(409), ack => zeropad3D_CP_2152_elements(975), clk => clk, reset =>reset);
    -- CP-element group 976:  transition  input  bypass 
    -- CP-element group 976: predecessors 
    -- CP-element group 976: 	409 
    -- CP-element group 976: successors 
    -- CP-element group 976: 	978 
    -- CP-element group 976:  members (2) 
      -- CP-element group 976: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2995/SplitProtocol/Sample/ra
      -- CP-element group 976: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2995/SplitProtocol/Sample/$exit
      -- 
    ra_12480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 976_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2995_inst_ack_0, ack => zeropad3D_CP_2152_elements(976)); -- 
    -- CP-element group 977:  transition  input  bypass 
    -- CP-element group 977: predecessors 
    -- CP-element group 977: 	409 
    -- CP-element group 977: successors 
    -- CP-element group 977: 	978 
    -- CP-element group 977:  members (2) 
      -- CP-element group 977: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2995/SplitProtocol/Update/ca
      -- CP-element group 977: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2995/SplitProtocol/Update/$exit
      -- 
    ca_12485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 977_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2995_inst_ack_1, ack => zeropad3D_CP_2152_elements(977)); -- 
    -- CP-element group 978:  join  transition  output  bypass 
    -- CP-element group 978: predecessors 
    -- CP-element group 978: 	976 
    -- CP-element group 978: 	977 
    -- CP-element group 978: successors 
    -- CP-element group 978: 	982 
    -- CP-element group 978:  members (5) 
      -- CP-element group 978: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_req
      -- CP-element group 978: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2995/SplitProtocol/$exit
      -- CP-element group 978: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2995/$exit
      -- CP-element group 978: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/$exit
      -- CP-element group 978: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2990/$exit
      -- 
    phi_stmt_2990_req_12486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2990_req_12486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(978), ack => phi_stmt_2990_req_1); -- 
    zeropad3D_cp_element_group_978: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_978"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(976) & zeropad3D_CP_2152_elements(977);
      gj_zeropad3D_cp_element_group_978 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(978), clk => clk, reset => reset); --
    end block;
    -- CP-element group 979:  transition  input  bypass 
    -- CP-element group 979: predecessors 
    -- CP-element group 979: 	409 
    -- CP-element group 979: successors 
    -- CP-element group 979: 	981 
    -- CP-element group 979:  members (2) 
      -- CP-element group 979: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_3001/SplitProtocol/Sample/ra
      -- CP-element group 979: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_3001/SplitProtocol/Sample/$exit
      -- 
    ra_12503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 979_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3001_inst_ack_0, ack => zeropad3D_CP_2152_elements(979)); -- 
    -- CP-element group 980:  transition  input  bypass 
    -- CP-element group 980: predecessors 
    -- CP-element group 980: 	409 
    -- CP-element group 980: successors 
    -- CP-element group 980: 	981 
    -- CP-element group 980:  members (2) 
      -- CP-element group 980: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_3001/SplitProtocol/Update/ca
      -- CP-element group 980: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_3001/SplitProtocol/Update/$exit
      -- 
    ca_12508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 980_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3001_inst_ack_1, ack => zeropad3D_CP_2152_elements(980)); -- 
    -- CP-element group 981:  join  transition  output  bypass 
    -- CP-element group 981: predecessors 
    -- CP-element group 981: 	979 
    -- CP-element group 981: 	980 
    -- CP-element group 981: successors 
    -- CP-element group 981: 	982 
    -- CP-element group 981:  members (5) 
      -- CP-element group 981: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_3001/$exit
      -- CP-element group 981: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/$exit
      -- CP-element group 981: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/$exit
      -- CP-element group 981: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_req
      -- CP-element group 981: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_3001/SplitProtocol/$exit
      -- 
    phi_stmt_2996_req_12509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2996_req_12509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(981), ack => phi_stmt_2996_req_1); -- 
    zeropad3D_cp_element_group_981: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_981"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(979) & zeropad3D_CP_2152_elements(980);
      gj_zeropad3D_cp_element_group_981 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(981), clk => clk, reset => reset); --
    end block;
    -- CP-element group 982:  join  transition  bypass 
    -- CP-element group 982: predecessors 
    -- CP-element group 982: 	975 
    -- CP-element group 982: 	978 
    -- CP-element group 982: 	981 
    -- CP-element group 982: successors 
    -- CP-element group 982: 	993 
    -- CP-element group 982:  members (1) 
      -- CP-element group 982: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_982: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_982"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(975) & zeropad3D_CP_2152_elements(978) & zeropad3D_CP_2152_elements(981);
      gj_zeropad3D_cp_element_group_982 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(982), clk => clk, reset => reset); --
    end block;
    -- CP-element group 983:  transition  input  bypass 
    -- CP-element group 983: predecessors 
    -- CP-element group 983: 	390 
    -- CP-element group 983: successors 
    -- CP-element group 983: 	985 
    -- CP-element group 983:  members (2) 
      -- CP-element group 983: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/type_cast_2986/SplitProtocol/Sample/$exit
      -- CP-element group 983: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/type_cast_2986/SplitProtocol/Sample/ra
      -- 
    ra_12529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 983_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2986_inst_ack_0, ack => zeropad3D_CP_2152_elements(983)); -- 
    -- CP-element group 984:  transition  input  bypass 
    -- CP-element group 984: predecessors 
    -- CP-element group 984: 	390 
    -- CP-element group 984: successors 
    -- CP-element group 984: 	985 
    -- CP-element group 984:  members (2) 
      -- CP-element group 984: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/type_cast_2986/SplitProtocol/Update/ca
      -- CP-element group 984: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/type_cast_2986/SplitProtocol/Update/$exit
      -- 
    ca_12534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 984_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2986_inst_ack_1, ack => zeropad3D_CP_2152_elements(984)); -- 
    -- CP-element group 985:  join  transition  output  bypass 
    -- CP-element group 985: predecessors 
    -- CP-element group 985: 	983 
    -- CP-element group 985: 	984 
    -- CP-element group 985: successors 
    -- CP-element group 985: 	992 
    -- CP-element group 985:  members (5) 
      -- CP-element group 985: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/type_cast_2986/$exit
      -- CP-element group 985: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/type_cast_2986/SplitProtocol/$exit
      -- CP-element group 985: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_sources/$exit
      -- CP-element group 985: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/$exit
      -- CP-element group 985: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2983/phi_stmt_2983_req
      -- 
    phi_stmt_2983_req_12535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2983_req_12535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(985), ack => phi_stmt_2983_req_0); -- 
    zeropad3D_cp_element_group_985: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_985"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(983) & zeropad3D_CP_2152_elements(984);
      gj_zeropad3D_cp_element_group_985 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(985), clk => clk, reset => reset); --
    end block;
    -- CP-element group 986:  transition  input  bypass 
    -- CP-element group 986: predecessors 
    -- CP-element group 986: 	390 
    -- CP-element group 986: successors 
    -- CP-element group 986: 	988 
    -- CP-element group 986:  members (2) 
      -- CP-element group 986: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/$exit
      -- CP-element group 986: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/ra
      -- 
    ra_12552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 986_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2993_inst_ack_0, ack => zeropad3D_CP_2152_elements(986)); -- 
    -- CP-element group 987:  transition  input  bypass 
    -- CP-element group 987: predecessors 
    -- CP-element group 987: 	390 
    -- CP-element group 987: successors 
    -- CP-element group 987: 	988 
    -- CP-element group 987:  members (2) 
      -- CP-element group 987: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/ca
      -- CP-element group 987: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/$exit
      -- 
    ca_12557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 987_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2993_inst_ack_1, ack => zeropad3D_CP_2152_elements(987)); -- 
    -- CP-element group 988:  join  transition  output  bypass 
    -- CP-element group 988: predecessors 
    -- CP-element group 988: 	986 
    -- CP-element group 988: 	987 
    -- CP-element group 988: successors 
    -- CP-element group 988: 	992 
    -- CP-element group 988:  members (5) 
      -- CP-element group 988: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/$exit
      -- CP-element group 988: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/$exit
      -- CP-element group 988: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/$exit
      -- CP-element group 988: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/$exit
      -- CP-element group 988: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2990/phi_stmt_2990_req
      -- 
    phi_stmt_2990_req_12558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2990_req_12558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(988), ack => phi_stmt_2990_req_0); -- 
    zeropad3D_cp_element_group_988: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_988"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(986) & zeropad3D_CP_2152_elements(987);
      gj_zeropad3D_cp_element_group_988 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(988), clk => clk, reset => reset); --
    end block;
    -- CP-element group 989:  transition  input  bypass 
    -- CP-element group 989: predecessors 
    -- CP-element group 989: 	390 
    -- CP-element group 989: successors 
    -- CP-element group 989: 	991 
    -- CP-element group 989:  members (2) 
      -- CP-element group 989: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_2999/SplitProtocol/Sample/ra
      -- CP-element group 989: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_2999/SplitProtocol/Sample/$exit
      -- 
    ra_12575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 989_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2999_inst_ack_0, ack => zeropad3D_CP_2152_elements(989)); -- 
    -- CP-element group 990:  transition  input  bypass 
    -- CP-element group 990: predecessors 
    -- CP-element group 990: 	390 
    -- CP-element group 990: successors 
    -- CP-element group 990: 	991 
    -- CP-element group 990:  members (2) 
      -- CP-element group 990: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_2999/SplitProtocol/Update/ca
      -- CP-element group 990: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_2999/SplitProtocol/Update/$exit
      -- 
    ca_12580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 990_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2999_inst_ack_1, ack => zeropad3D_CP_2152_elements(990)); -- 
    -- CP-element group 991:  join  transition  output  bypass 
    -- CP-element group 991: predecessors 
    -- CP-element group 991: 	989 
    -- CP-element group 991: 	990 
    -- CP-element group 991: successors 
    -- CP-element group 991: 	992 
    -- CP-element group 991:  members (5) 
      -- CP-element group 991: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_req
      -- CP-element group 991: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_2999/SplitProtocol/$exit
      -- CP-element group 991: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/type_cast_2999/$exit
      -- CP-element group 991: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/phi_stmt_2996_sources/$exit
      -- CP-element group 991: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2996/$exit
      -- 
    phi_stmt_2996_req_12581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2996_req_12581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(991), ack => phi_stmt_2996_req_0); -- 
    zeropad3D_cp_element_group_991: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_991"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(989) & zeropad3D_CP_2152_elements(990);
      gj_zeropad3D_cp_element_group_991 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(991), clk => clk, reset => reset); --
    end block;
    -- CP-element group 992:  join  transition  bypass 
    -- CP-element group 992: predecessors 
    -- CP-element group 992: 	985 
    -- CP-element group 992: 	988 
    -- CP-element group 992: 	991 
    -- CP-element group 992: successors 
    -- CP-element group 992: 	993 
    -- CP-element group 992:  members (1) 
      -- CP-element group 992: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_992: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_992"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(985) & zeropad3D_CP_2152_elements(988) & zeropad3D_CP_2152_elements(991);
      gj_zeropad3D_cp_element_group_992 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(992), clk => clk, reset => reset); --
    end block;
    -- CP-element group 993:  merge  fork  transition  place  bypass 
    -- CP-element group 993: predecessors 
    -- CP-element group 993: 	982 
    -- CP-element group 993: 	992 
    -- CP-element group 993: successors 
    -- CP-element group 993: 	994 
    -- CP-element group 993: 	995 
    -- CP-element group 993: 	996 
    -- CP-element group 993:  members (2) 
      -- CP-element group 993: 	 branch_block_stmt_714/merge_stmt_2982_PhiReqMerge
      -- CP-element group 993: 	 branch_block_stmt_714/merge_stmt_2982_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(993) <= OrReduce(zeropad3D_CP_2152_elements(982) & zeropad3D_CP_2152_elements(992));
    -- CP-element group 994:  transition  input  bypass 
    -- CP-element group 994: predecessors 
    -- CP-element group 994: 	993 
    -- CP-element group 994: successors 
    -- CP-element group 994: 	997 
    -- CP-element group 994:  members (1) 
      -- CP-element group 994: 	 branch_block_stmt_714/merge_stmt_2982_PhiAck/phi_stmt_2983_ack
      -- 
    phi_stmt_2983_ack_12586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 994_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2983_ack_0, ack => zeropad3D_CP_2152_elements(994)); -- 
    -- CP-element group 995:  transition  input  bypass 
    -- CP-element group 995: predecessors 
    -- CP-element group 995: 	993 
    -- CP-element group 995: successors 
    -- CP-element group 995: 	997 
    -- CP-element group 995:  members (1) 
      -- CP-element group 995: 	 branch_block_stmt_714/merge_stmt_2982_PhiAck/phi_stmt_2990_ack
      -- 
    phi_stmt_2990_ack_12587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 995_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2990_ack_0, ack => zeropad3D_CP_2152_elements(995)); -- 
    -- CP-element group 996:  transition  input  bypass 
    -- CP-element group 996: predecessors 
    -- CP-element group 996: 	993 
    -- CP-element group 996: successors 
    -- CP-element group 996: 	997 
    -- CP-element group 996:  members (1) 
      -- CP-element group 996: 	 branch_block_stmt_714/merge_stmt_2982_PhiAck/phi_stmt_2996_ack
      -- 
    phi_stmt_2996_ack_12588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 996_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2996_ack_0, ack => zeropad3D_CP_2152_elements(996)); -- 
    -- CP-element group 997:  join  transition  bypass 
    -- CP-element group 997: predecessors 
    -- CP-element group 997: 	994 
    -- CP-element group 997: 	995 
    -- CP-element group 997: 	996 
    -- CP-element group 997: successors 
    -- CP-element group 997: 	4 
    -- CP-element group 997:  members (1) 
      -- CP-element group 997: 	 branch_block_stmt_714/merge_stmt_2982_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_997: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_997"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(994) & zeropad3D_CP_2152_elements(995) & zeropad3D_CP_2152_elements(996);
      gj_zeropad3D_cp_element_group_997 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(997), clk => clk, reset => reset); --
    end block;
    -- CP-element group 998:  transition  input  bypass 
    -- CP-element group 998: predecessors 
    -- CP-element group 998: 	408 
    -- CP-element group 998: successors 
    -- CP-element group 998: 	1000 
    -- CP-element group 998:  members (2) 
      -- CP-element group 998: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3008/SplitProtocol/Sample/ra
      -- CP-element group 998: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3008/SplitProtocol/Sample/$exit
      -- 
    ra_12608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 998_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3008_inst_ack_0, ack => zeropad3D_CP_2152_elements(998)); -- 
    -- CP-element group 999:  transition  input  bypass 
    -- CP-element group 999: predecessors 
    -- CP-element group 999: 	408 
    -- CP-element group 999: successors 
    -- CP-element group 999: 	1000 
    -- CP-element group 999:  members (2) 
      -- CP-element group 999: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3008/SplitProtocol/Update/ca
      -- CP-element group 999: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3008/SplitProtocol/Update/$exit
      -- 
    ca_12613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 999_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3008_inst_ack_1, ack => zeropad3D_CP_2152_elements(999)); -- 
    -- CP-element group 1000:  join  transition  output  bypass 
    -- CP-element group 1000: predecessors 
    -- CP-element group 1000: 	998 
    -- CP-element group 1000: 	999 
    -- CP-element group 1000: successors 
    -- CP-element group 1000: 	1004 
    -- CP-element group 1000:  members (5) 
      -- CP-element group 1000: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_req
      -- CP-element group 1000: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3008/SplitProtocol/$exit
      -- CP-element group 1000: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3008/$exit
      -- CP-element group 1000: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/$exit
      -- CP-element group 1000: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3005/$exit
      -- 
    phi_stmt_3005_req_12614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3005_req_12614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1000), ack => phi_stmt_3005_req_0); -- 
    zeropad3D_cp_element_group_1000: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1000"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(998) & zeropad3D_CP_2152_elements(999);
      gj_zeropad3D_cp_element_group_1000 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1000), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1001:  transition  input  bypass 
    -- CP-element group 1001: predecessors 
    -- CP-element group 1001: 	408 
    -- CP-element group 1001: successors 
    -- CP-element group 1001: 	1003 
    -- CP-element group 1001:  members (2) 
      -- CP-element group 1001: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/type_cast_3012/SplitProtocol/Sample/$exit
      -- CP-element group 1001: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/type_cast_3012/SplitProtocol/Sample/ra
      -- 
    ra_12631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1001_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3012_inst_ack_0, ack => zeropad3D_CP_2152_elements(1001)); -- 
    -- CP-element group 1002:  transition  input  bypass 
    -- CP-element group 1002: predecessors 
    -- CP-element group 1002: 	408 
    -- CP-element group 1002: successors 
    -- CP-element group 1002: 	1003 
    -- CP-element group 1002:  members (2) 
      -- CP-element group 1002: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/type_cast_3012/SplitProtocol/Update/$exit
      -- CP-element group 1002: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/type_cast_3012/SplitProtocol/Update/ca
      -- 
    ca_12636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1002_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3012_inst_ack_1, ack => zeropad3D_CP_2152_elements(1002)); -- 
    -- CP-element group 1003:  join  transition  output  bypass 
    -- CP-element group 1003: predecessors 
    -- CP-element group 1003: 	1001 
    -- CP-element group 1003: 	1002 
    -- CP-element group 1003: successors 
    -- CP-element group 1003: 	1004 
    -- CP-element group 1003:  members (5) 
      -- CP-element group 1003: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_req
      -- CP-element group 1003: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/$exit
      -- CP-element group 1003: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/type_cast_3012/SplitProtocol/$exit
      -- CP-element group 1003: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/type_cast_3012/$exit
      -- CP-element group 1003: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/phi_stmt_3009/phi_stmt_3009_sources/$exit
      -- 
    phi_stmt_3009_req_12637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3009_req_12637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1003), ack => phi_stmt_3009_req_0); -- 
    zeropad3D_cp_element_group_1003: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1003"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1001) & zeropad3D_CP_2152_elements(1002);
      gj_zeropad3D_cp_element_group_1003 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1003), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1004:  join  fork  transition  place  bypass 
    -- CP-element group 1004: predecessors 
    -- CP-element group 1004: 	1000 
    -- CP-element group 1004: 	1003 
    -- CP-element group 1004: successors 
    -- CP-element group 1004: 	1005 
    -- CP-element group 1004: 	1006 
    -- CP-element group 1004:  members (3) 
      -- CP-element group 1004: 	 branch_block_stmt_714/merge_stmt_3004_PhiReqMerge
      -- CP-element group 1004: 	 branch_block_stmt_714/merge_stmt_3004_PhiAck/$entry
      -- CP-element group 1004: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1004: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1004"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1000) & zeropad3D_CP_2152_elements(1003);
      gj_zeropad3D_cp_element_group_1004 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1004), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1005:  transition  input  bypass 
    -- CP-element group 1005: predecessors 
    -- CP-element group 1005: 	1004 
    -- CP-element group 1005: successors 
    -- CP-element group 1005: 	1007 
    -- CP-element group 1005:  members (1) 
      -- CP-element group 1005: 	 branch_block_stmt_714/merge_stmt_3004_PhiAck/phi_stmt_3005_ack
      -- 
    phi_stmt_3005_ack_12642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1005_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3005_ack_0, ack => zeropad3D_CP_2152_elements(1005)); -- 
    -- CP-element group 1006:  transition  input  bypass 
    -- CP-element group 1006: predecessors 
    -- CP-element group 1006: 	1004 
    -- CP-element group 1006: successors 
    -- CP-element group 1006: 	1007 
    -- CP-element group 1006:  members (1) 
      -- CP-element group 1006: 	 branch_block_stmt_714/merge_stmt_3004_PhiAck/phi_stmt_3009_ack
      -- 
    phi_stmt_3009_ack_12643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1006_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3009_ack_0, ack => zeropad3D_CP_2152_elements(1006)); -- 
    -- CP-element group 1007:  join  fork  transition  place  output  bypass 
    -- CP-element group 1007: predecessors 
    -- CP-element group 1007: 	1005 
    -- CP-element group 1007: 	1006 
    -- CP-element group 1007: successors 
    -- CP-element group 1007: 	410 
    -- CP-element group 1007: 	411 
    -- CP-element group 1007: 	412 
    -- CP-element group 1007: 	413 
    -- CP-element group 1007: 	414 
    -- CP-element group 1007: 	415 
    -- CP-element group 1007: 	416 
    -- CP-element group 1007: 	417 
    -- CP-element group 1007: 	418 
    -- CP-element group 1007: 	419 
    -- CP-element group 1007: 	421 
    -- CP-element group 1007: 	423 
    -- CP-element group 1007:  members (92) 
      -- CP-element group 1007: 	 branch_block_stmt_714/merge_stmt_3004__exit__
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137__entry__
      -- CP-element group 1007: 	 branch_block_stmt_714/merge_stmt_3004_PhiAck/$exit
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3016_sample_start_
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3016_update_start_
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3016_Sample/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3016_Sample/rr
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3016_Update/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3016_Update/cr
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_sample_start_
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_update_start_
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_word_address_calculated
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_root_address_calculated
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Sample/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Sample/word_access_start/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Sample/word_access_start/word_0/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Sample/word_access_start/word_0/rr
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Update/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Update/word_access_complete/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Update/word_access_complete/word_0/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_pad_3025_Update/word_access_complete/word_0/cr
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_sample_start_
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_update_start_
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_word_address_calculated
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_root_address_calculated
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Sample/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Sample/word_access_start/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Sample/word_access_start/word_0/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Sample/word_access_start/word_0/rr
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Update/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Update/word_access_complete/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Update/word_access_complete/word_0/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/LOAD_depth_high_3028_Update/word_access_complete/word_0/cr
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_sample_start_
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_update_start_
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_base_address_calculated
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_word_address_calculated
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_root_address_calculated
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_base_address_resized
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_base_addr_resize/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_base_addr_resize/$exit
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_base_addr_resize/base_resize_req
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_base_addr_resize/base_resize_ack
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_base_plus_offset/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_base_plus_offset/$exit
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_base_plus_offset/sum_rename_req
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_base_plus_offset/sum_rename_ack
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_word_addrgen/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_word_addrgen/$exit
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_word_addrgen/root_register_req
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_word_addrgen/root_register_ack
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Sample/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Sample/word_access_start/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Sample/word_access_start/word_0/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Sample/word_access_start/word_0/rr
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Update/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Update/word_access_complete/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Update/word_access_complete/word_0/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3040_Update/word_access_complete/word_0/cr
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_sample_start_
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_update_start_
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_base_address_calculated
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_word_address_calculated
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_root_address_calculated
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_base_address_resized
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_base_addr_resize/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_base_addr_resize/$exit
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_base_addr_resize/base_resize_req
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_base_addr_resize/base_resize_ack
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_base_plus_offset/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_base_plus_offset/$exit
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_base_plus_offset/sum_rename_req
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_base_plus_offset/sum_rename_ack
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_word_addrgen/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_word_addrgen/$exit
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_word_addrgen/root_register_req
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_word_addrgen/root_register_ack
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Sample/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Sample/word_access_start/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Sample/word_access_start/word_0/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Sample/word_access_start/word_0/rr
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Update/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Update/word_access_complete/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Update/word_access_complete/word_0/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/ptr_deref_3052_Update/word_access_complete/word_0/cr
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3056_update_start_
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3056_Update/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3056_Update/cr
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3095_update_start_
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3095_Update/$entry
      -- CP-element group 1007: 	 branch_block_stmt_714/assign_stmt_3017_to_assign_stmt_3137/type_cast_3095_Update/cr
      -- 
    rr_6953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1007), ack => type_cast_3016_inst_req_0); -- 
    cr_6958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1007), ack => type_cast_3016_inst_req_1); -- 
    rr_6975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1007), ack => LOAD_pad_3025_load_0_req_0); -- 
    cr_6986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1007), ack => LOAD_pad_3025_load_0_req_1); -- 
    rr_7008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1007), ack => LOAD_depth_high_3028_load_0_req_0); -- 
    cr_7019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1007), ack => LOAD_depth_high_3028_load_0_req_1); -- 
    rr_7058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1007), ack => ptr_deref_3040_load_0_req_0); -- 
    cr_7069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1007), ack => ptr_deref_3040_load_0_req_1); -- 
    rr_7108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1007), ack => ptr_deref_3052_load_0_req_0); -- 
    cr_7119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1007), ack => ptr_deref_3052_load_0_req_1); -- 
    cr_7138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1007), ack => type_cast_3056_inst_req_1); -- 
    cr_7152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1007), ack => type_cast_3095_inst_req_1); -- 
    zeropad3D_cp_element_group_1007: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1007"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1005) & zeropad3D_CP_2152_elements(1006);
      gj_zeropad3D_cp_element_group_1007 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1007), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1008:  transition  input  bypass 
    -- CP-element group 1008: predecessors 
    -- CP-element group 1008: 	5 
    -- CP-element group 1008: successors 
    -- CP-element group 1008: 	1010 
    -- CP-element group 1008:  members (2) 
      -- CP-element group 1008: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/type_cast_3156/SplitProtocol/Sample/ra
      -- CP-element group 1008: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/type_cast_3156/SplitProtocol/Sample/$exit
      -- 
    ra_12663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1008_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3156_inst_ack_0, ack => zeropad3D_CP_2152_elements(1008)); -- 
    -- CP-element group 1009:  transition  input  bypass 
    -- CP-element group 1009: predecessors 
    -- CP-element group 1009: 	5 
    -- CP-element group 1009: successors 
    -- CP-element group 1009: 	1010 
    -- CP-element group 1009:  members (2) 
      -- CP-element group 1009: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/type_cast_3156/SplitProtocol/Update/ca
      -- CP-element group 1009: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/type_cast_3156/SplitProtocol/Update/$exit
      -- 
    ca_12668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1009_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3156_inst_ack_1, ack => zeropad3D_CP_2152_elements(1009)); -- 
    -- CP-element group 1010:  join  transition  output  bypass 
    -- CP-element group 1010: predecessors 
    -- CP-element group 1010: 	1008 
    -- CP-element group 1010: 	1009 
    -- CP-element group 1010: successors 
    -- CP-element group 1010: 	1017 
    -- CP-element group 1010:  members (5) 
      -- CP-element group 1010: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/type_cast_3156/$exit
      -- CP-element group 1010: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_req
      -- CP-element group 1010: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/$exit
      -- CP-element group 1010: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/$exit
      -- CP-element group 1010: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/type_cast_3156/SplitProtocol/$exit
      -- 
    phi_stmt_3153_req_12669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3153_req_12669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1010), ack => phi_stmt_3153_req_0); -- 
    zeropad3D_cp_element_group_1010: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1010"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1008) & zeropad3D_CP_2152_elements(1009);
      gj_zeropad3D_cp_element_group_1010 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1010), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1011:  transition  input  bypass 
    -- CP-element group 1011: predecessors 
    -- CP-element group 1011: 	5 
    -- CP-element group 1011: successors 
    -- CP-element group 1011: 	1013 
    -- CP-element group 1011:  members (2) 
      -- CP-element group 1011: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3150/SplitProtocol/Sample/ra
      -- CP-element group 1011: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3150/SplitProtocol/Sample/$exit
      -- 
    ra_12686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1011_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3150_inst_ack_0, ack => zeropad3D_CP_2152_elements(1011)); -- 
    -- CP-element group 1012:  transition  input  bypass 
    -- CP-element group 1012: predecessors 
    -- CP-element group 1012: 	5 
    -- CP-element group 1012: successors 
    -- CP-element group 1012: 	1013 
    -- CP-element group 1012:  members (2) 
      -- CP-element group 1012: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3150/SplitProtocol/Update/ca
      -- CP-element group 1012: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3150/SplitProtocol/Update/$exit
      -- 
    ca_12691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1012_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3150_inst_ack_1, ack => zeropad3D_CP_2152_elements(1012)); -- 
    -- CP-element group 1013:  join  transition  output  bypass 
    -- CP-element group 1013: predecessors 
    -- CP-element group 1013: 	1011 
    -- CP-element group 1013: 	1012 
    -- CP-element group 1013: successors 
    -- CP-element group 1013: 	1017 
    -- CP-element group 1013:  members (5) 
      -- CP-element group 1013: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_req
      -- CP-element group 1013: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3150/SplitProtocol/$exit
      -- CP-element group 1013: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3150/$exit
      -- CP-element group 1013: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/$exit
      -- CP-element group 1013: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3147/$exit
      -- 
    phi_stmt_3147_req_12692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3147_req_12692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1013), ack => phi_stmt_3147_req_0); -- 
    zeropad3D_cp_element_group_1013: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1013"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1011) & zeropad3D_CP_2152_elements(1012);
      gj_zeropad3D_cp_element_group_1013 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1013), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1014:  transition  input  bypass 
    -- CP-element group 1014: predecessors 
    -- CP-element group 1014: 	5 
    -- CP-element group 1014: successors 
    -- CP-element group 1014: 	1016 
    -- CP-element group 1014:  members (2) 
      -- CP-element group 1014: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/type_cast_3146/SplitProtocol/Sample/ra
      -- CP-element group 1014: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/type_cast_3146/SplitProtocol/Sample/$exit
      -- 
    ra_12709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1014_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3146_inst_ack_0, ack => zeropad3D_CP_2152_elements(1014)); -- 
    -- CP-element group 1015:  transition  input  bypass 
    -- CP-element group 1015: predecessors 
    -- CP-element group 1015: 	5 
    -- CP-element group 1015: successors 
    -- CP-element group 1015: 	1016 
    -- CP-element group 1015:  members (2) 
      -- CP-element group 1015: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/type_cast_3146/SplitProtocol/Update/ca
      -- CP-element group 1015: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/type_cast_3146/SplitProtocol/Update/$exit
      -- 
    ca_12714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1015_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3146_inst_ack_1, ack => zeropad3D_CP_2152_elements(1015)); -- 
    -- CP-element group 1016:  join  transition  output  bypass 
    -- CP-element group 1016: predecessors 
    -- CP-element group 1016: 	1014 
    -- CP-element group 1016: 	1015 
    -- CP-element group 1016: successors 
    -- CP-element group 1016: 	1017 
    -- CP-element group 1016:  members (5) 
      -- CP-element group 1016: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/$exit
      -- CP-element group 1016: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/type_cast_3146/$exit
      -- CP-element group 1016: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/$exit
      -- CP-element group 1016: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/type_cast_3146/SplitProtocol/$exit
      -- CP-element group 1016: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_req
      -- 
    phi_stmt_3140_req_12715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3140_req_12715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1016), ack => phi_stmt_3140_req_1); -- 
    zeropad3D_cp_element_group_1016: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1016"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1014) & zeropad3D_CP_2152_elements(1015);
      gj_zeropad3D_cp_element_group_1016 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1016), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1017:  join  transition  bypass 
    -- CP-element group 1017: predecessors 
    -- CP-element group 1017: 	1010 
    -- CP-element group 1017: 	1013 
    -- CP-element group 1017: 	1016 
    -- CP-element group 1017: successors 
    -- CP-element group 1017: 	1024 
    -- CP-element group 1017:  members (1) 
      -- CP-element group 1017: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1017: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1017"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1010) & zeropad3D_CP_2152_elements(1013) & zeropad3D_CP_2152_elements(1016);
      gj_zeropad3D_cp_element_group_1017 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1017), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1018:  transition  output  delay-element  bypass 
    -- CP-element group 1018: predecessors 
    -- CP-element group 1018: 	424 
    -- CP-element group 1018: successors 
    -- CP-element group 1018: 	1023 
    -- CP-element group 1018:  members (4) 
      -- CP-element group 1018: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_req
      -- CP-element group 1018: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/type_cast_3159_konst_delay_trans
      -- CP-element group 1018: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3153/phi_stmt_3153_sources/$exit
      -- CP-element group 1018: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3153/$exit
      -- 
    phi_stmt_3153_req_12726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3153_req_12726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1018), ack => phi_stmt_3153_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(1018) is a control-delay.
    cp_element_1018_delay: control_delay_element  generic map(name => " 1018_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(424), ack => zeropad3D_CP_2152_elements(1018), clk => clk, reset =>reset);
    -- CP-element group 1019:  transition  input  bypass 
    -- CP-element group 1019: predecessors 
    -- CP-element group 1019: 	424 
    -- CP-element group 1019: successors 
    -- CP-element group 1019: 	1021 
    -- CP-element group 1019:  members (2) 
      -- CP-element group 1019: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3152/SplitProtocol/Sample/ra
      -- CP-element group 1019: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3152/SplitProtocol/Sample/$exit
      -- 
    ra_12743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1019_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3152_inst_ack_0, ack => zeropad3D_CP_2152_elements(1019)); -- 
    -- CP-element group 1020:  transition  input  bypass 
    -- CP-element group 1020: predecessors 
    -- CP-element group 1020: 	424 
    -- CP-element group 1020: successors 
    -- CP-element group 1020: 	1021 
    -- CP-element group 1020:  members (2) 
      -- CP-element group 1020: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3152/SplitProtocol/Update/ca
      -- CP-element group 1020: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3152/SplitProtocol/Update/$exit
      -- 
    ca_12748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1020_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3152_inst_ack_1, ack => zeropad3D_CP_2152_elements(1020)); -- 
    -- CP-element group 1021:  join  transition  output  bypass 
    -- CP-element group 1021: predecessors 
    -- CP-element group 1021: 	1019 
    -- CP-element group 1021: 	1020 
    -- CP-element group 1021: successors 
    -- CP-element group 1021: 	1023 
    -- CP-element group 1021:  members (5) 
      -- CP-element group 1021: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/$exit
      -- CP-element group 1021: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/$exit
      -- CP-element group 1021: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_req
      -- CP-element group 1021: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3152/SplitProtocol/$exit
      -- CP-element group 1021: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3147/phi_stmt_3147_sources/type_cast_3152/$exit
      -- 
    phi_stmt_3147_req_12749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3147_req_12749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1021), ack => phi_stmt_3147_req_1); -- 
    zeropad3D_cp_element_group_1021: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1021"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1019) & zeropad3D_CP_2152_elements(1020);
      gj_zeropad3D_cp_element_group_1021 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1021), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1022:  transition  output  delay-element  bypass 
    -- CP-element group 1022: predecessors 
    -- CP-element group 1022: 	424 
    -- CP-element group 1022: successors 
    -- CP-element group 1022: 	1023 
    -- CP-element group 1022:  members (4) 
      -- CP-element group 1022: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_req
      -- CP-element group 1022: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/type_cast_3144_konst_delay_trans
      -- CP-element group 1022: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3140/phi_stmt_3140_sources/$exit
      -- CP-element group 1022: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3140/$exit
      -- 
    phi_stmt_3140_req_12757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3140_req_12757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1022), ack => phi_stmt_3140_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(1022) is a control-delay.
    cp_element_1022_delay: control_delay_element  generic map(name => " 1022_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(424), ack => zeropad3D_CP_2152_elements(1022), clk => clk, reset =>reset);
    -- CP-element group 1023:  join  transition  bypass 
    -- CP-element group 1023: predecessors 
    -- CP-element group 1023: 	1018 
    -- CP-element group 1023: 	1021 
    -- CP-element group 1023: 	1022 
    -- CP-element group 1023: successors 
    -- CP-element group 1023: 	1024 
    -- CP-element group 1023:  members (1) 
      -- CP-element group 1023: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1023: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1023"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1018) & zeropad3D_CP_2152_elements(1021) & zeropad3D_CP_2152_elements(1022);
      gj_zeropad3D_cp_element_group_1023 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1023), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1024:  merge  fork  transition  place  bypass 
    -- CP-element group 1024: predecessors 
    -- CP-element group 1024: 	1017 
    -- CP-element group 1024: 	1023 
    -- CP-element group 1024: successors 
    -- CP-element group 1024: 	1025 
    -- CP-element group 1024: 	1026 
    -- CP-element group 1024: 	1027 
    -- CP-element group 1024:  members (2) 
      -- CP-element group 1024: 	 branch_block_stmt_714/merge_stmt_3139_PhiAck/$entry
      -- CP-element group 1024: 	 branch_block_stmt_714/merge_stmt_3139_PhiReqMerge
      -- 
    zeropad3D_CP_2152_elements(1024) <= OrReduce(zeropad3D_CP_2152_elements(1017) & zeropad3D_CP_2152_elements(1023));
    -- CP-element group 1025:  transition  input  bypass 
    -- CP-element group 1025: predecessors 
    -- CP-element group 1025: 	1024 
    -- CP-element group 1025: successors 
    -- CP-element group 1025: 	1028 
    -- CP-element group 1025:  members (1) 
      -- CP-element group 1025: 	 branch_block_stmt_714/merge_stmt_3139_PhiAck/phi_stmt_3140_ack
      -- 
    phi_stmt_3140_ack_12762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1025_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3140_ack_0, ack => zeropad3D_CP_2152_elements(1025)); -- 
    -- CP-element group 1026:  transition  input  bypass 
    -- CP-element group 1026: predecessors 
    -- CP-element group 1026: 	1024 
    -- CP-element group 1026: successors 
    -- CP-element group 1026: 	1028 
    -- CP-element group 1026:  members (1) 
      -- CP-element group 1026: 	 branch_block_stmt_714/merge_stmt_3139_PhiAck/phi_stmt_3147_ack
      -- 
    phi_stmt_3147_ack_12763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1026_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3147_ack_0, ack => zeropad3D_CP_2152_elements(1026)); -- 
    -- CP-element group 1027:  transition  input  bypass 
    -- CP-element group 1027: predecessors 
    -- CP-element group 1027: 	1024 
    -- CP-element group 1027: successors 
    -- CP-element group 1027: 	1028 
    -- CP-element group 1027:  members (1) 
      -- CP-element group 1027: 	 branch_block_stmt_714/merge_stmt_3139_PhiAck/phi_stmt_3153_ack
      -- 
    phi_stmt_3153_ack_12764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1027_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3153_ack_0, ack => zeropad3D_CP_2152_elements(1027)); -- 
    -- CP-element group 1028:  join  fork  transition  place  output  bypass 
    -- CP-element group 1028: predecessors 
    -- CP-element group 1028: 	1025 
    -- CP-element group 1028: 	1026 
    -- CP-element group 1028: 	1027 
    -- CP-element group 1028: successors 
    -- CP-element group 1028: 	425 
    -- CP-element group 1028: 	426 
    -- CP-element group 1028:  members (10) 
      -- CP-element group 1028: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172__entry__
      -- CP-element group 1028: 	 branch_block_stmt_714/merge_stmt_3139__exit__
      -- CP-element group 1028: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/$entry
      -- CP-element group 1028: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/type_cast_3164_sample_start_
      -- CP-element group 1028: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/type_cast_3164_update_start_
      -- CP-element group 1028: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/type_cast_3164_Sample/$entry
      -- CP-element group 1028: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/type_cast_3164_Sample/rr
      -- CP-element group 1028: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/type_cast_3164_Update/$entry
      -- CP-element group 1028: 	 branch_block_stmt_714/assign_stmt_3165_to_assign_stmt_3172/type_cast_3164_Update/cr
      -- CP-element group 1028: 	 branch_block_stmt_714/merge_stmt_3139_PhiAck/$exit
      -- 
    rr_7164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1028), ack => type_cast_3164_inst_req_0); -- 
    cr_7169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1028), ack => type_cast_3164_inst_req_1); -- 
    zeropad3D_cp_element_group_1028: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1028"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1025) & zeropad3D_CP_2152_elements(1026) & zeropad3D_CP_2152_elements(1027);
      gj_zeropad3D_cp_element_group_1028 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1028), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1029:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1029: predecessors 
    -- CP-element group 1029: 	427 
    -- CP-element group 1029: 	434 
    -- CP-element group 1029: 	437 
    -- CP-element group 1029: 	444 
    -- CP-element group 1029: successors 
    -- CP-element group 1029: 	445 
    -- CP-element group 1029: 	446 
    -- CP-element group 1029: 	447 
    -- CP-element group 1029: 	448 
    -- CP-element group 1029: 	451 
    -- CP-element group 1029: 	453 
    -- CP-element group 1029: 	455 
    -- CP-element group 1029: 	457 
    -- CP-element group 1029:  members (33) 
      -- CP-element group 1029: 	 branch_block_stmt_714/merge_stmt_3268__exit__
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324__entry__
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/$entry
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3272_sample_start_
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3272_update_start_
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3272_Sample/$entry
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3272_Sample/rr
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3272_Update/$entry
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3272_Update/cr
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3277_sample_start_
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3277_update_start_
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3277_Sample/$entry
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3277_Sample/rr
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3277_Update/$entry
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3277_Update/cr
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3311_update_start_
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3311_Update/$entry
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/type_cast_3311_Update/cr
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/addr_of_3318_update_start_
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_final_index_sum_regn_update_start
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_final_index_sum_regn_Update/$entry
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/array_obj_ref_3317_final_index_sum_regn_Update/req
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/addr_of_3318_complete/$entry
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/addr_of_3318_complete/req
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_update_start_
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Update/$entry
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Update/word_access_complete/$entry
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Update/word_access_complete/word_0/$entry
      -- CP-element group 1029: 	 branch_block_stmt_714/assign_stmt_3273_to_assign_stmt_3324/ptr_deref_3321_Update/word_access_complete/word_0/cr
      -- CP-element group 1029: 	 branch_block_stmt_714/merge_stmt_3268_PhiReqMerge
      -- CP-element group 1029: 	 branch_block_stmt_714/merge_stmt_3268_PhiAck/$entry
      -- CP-element group 1029: 	 branch_block_stmt_714/merge_stmt_3268_PhiAck/$exit
      -- CP-element group 1029: 	 branch_block_stmt_714/merge_stmt_3268_PhiAck/dummy
      -- 
    rr_7374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1029), ack => type_cast_3272_inst_req_0); -- 
    cr_7379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1029), ack => type_cast_3272_inst_req_1); -- 
    rr_7388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1029), ack => type_cast_3277_inst_req_0); -- 
    cr_7393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1029), ack => type_cast_3277_inst_req_1); -- 
    cr_7407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1029), ack => type_cast_3311_inst_req_1); -- 
    req_7438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1029), ack => array_obj_ref_3317_index_offset_req_1); -- 
    req_7453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1029), ack => addr_of_3318_final_reg_req_1); -- 
    cr_7503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1029), ack => ptr_deref_3321_store_0_req_1); -- 
    zeropad3D_CP_2152_elements(1029) <= OrReduce(zeropad3D_CP_2152_elements(427) & zeropad3D_CP_2152_elements(434) & zeropad3D_CP_2152_elements(437) & zeropad3D_CP_2152_elements(444));
    -- CP-element group 1030:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1030: predecessors 
    -- CP-element group 1030: 	458 
    -- CP-element group 1030: 	478 
    -- CP-element group 1030: successors 
    -- CP-element group 1030: 	479 
    -- CP-element group 1030: 	480 
    -- CP-element group 1030:  members (13) 
      -- CP-element group 1030: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451__entry__
      -- CP-element group 1030: 	 branch_block_stmt_714/merge_stmt_3433__exit__
      -- CP-element group 1030: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/type_cast_3437_update_start_
      -- CP-element group 1030: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/type_cast_3437_Sample/$entry
      -- CP-element group 1030: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/type_cast_3437_Sample/rr
      -- CP-element group 1030: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/type_cast_3437_Update/$entry
      -- CP-element group 1030: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/type_cast_3437_sample_start_
      -- CP-element group 1030: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/$entry
      -- CP-element group 1030: 	 branch_block_stmt_714/assign_stmt_3438_to_assign_stmt_3451/type_cast_3437_Update/cr
      -- CP-element group 1030: 	 branch_block_stmt_714/merge_stmt_3433_PhiReqMerge
      -- CP-element group 1030: 	 branch_block_stmt_714/merge_stmt_3433_PhiAck/$entry
      -- CP-element group 1030: 	 branch_block_stmt_714/merge_stmt_3433_PhiAck/$exit
      -- CP-element group 1030: 	 branch_block_stmt_714/merge_stmt_3433_PhiAck/dummy
      -- 
    rr_7752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1030), ack => type_cast_3437_inst_req_0); -- 
    cr_7757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1030), ack => type_cast_3437_inst_req_1); -- 
    zeropad3D_CP_2152_elements(1030) <= OrReduce(zeropad3D_CP_2152_elements(458) & zeropad3D_CP_2152_elements(478));
    -- CP-element group 1031:  transition  output  delay-element  bypass 
    -- CP-element group 1031: predecessors 
    -- CP-element group 1031: 	500 
    -- CP-element group 1031: successors 
    -- CP-element group 1031: 	1038 
    -- CP-element group 1031:  members (4) 
      -- CP-element group 1031: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3558/$exit
      -- CP-element group 1031: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/$exit
      -- CP-element group 1031: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/type_cast_3564_konst_delay_trans
      -- CP-element group 1031: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_req
      -- 
    phi_stmt_3558_req_12875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3558_req_12875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1031), ack => phi_stmt_3558_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(1031) is a control-delay.
    cp_element_1031_delay: control_delay_element  generic map(name => " 1031_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(500), ack => zeropad3D_CP_2152_elements(1031), clk => clk, reset =>reset);
    -- CP-element group 1032:  transition  input  bypass 
    -- CP-element group 1032: predecessors 
    -- CP-element group 1032: 	500 
    -- CP-element group 1032: successors 
    -- CP-element group 1032: 	1034 
    -- CP-element group 1032:  members (2) 
      -- CP-element group 1032: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3570/SplitProtocol/Sample/$exit
      -- CP-element group 1032: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3570/SplitProtocol/Sample/ra
      -- 
    ra_12892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1032_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3570_inst_ack_0, ack => zeropad3D_CP_2152_elements(1032)); -- 
    -- CP-element group 1033:  transition  input  bypass 
    -- CP-element group 1033: predecessors 
    -- CP-element group 1033: 	500 
    -- CP-element group 1033: successors 
    -- CP-element group 1033: 	1034 
    -- CP-element group 1033:  members (2) 
      -- CP-element group 1033: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3570/SplitProtocol/Update/$exit
      -- CP-element group 1033: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3570/SplitProtocol/Update/ca
      -- 
    ca_12897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1033_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3570_inst_ack_1, ack => zeropad3D_CP_2152_elements(1033)); -- 
    -- CP-element group 1034:  join  transition  output  bypass 
    -- CP-element group 1034: predecessors 
    -- CP-element group 1034: 	1032 
    -- CP-element group 1034: 	1033 
    -- CP-element group 1034: successors 
    -- CP-element group 1034: 	1038 
    -- CP-element group 1034:  members (5) 
      -- CP-element group 1034: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/$exit
      -- CP-element group 1034: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/$exit
      -- CP-element group 1034: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3570/$exit
      -- CP-element group 1034: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3570/SplitProtocol/$exit
      -- CP-element group 1034: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_req
      -- 
    phi_stmt_3565_req_12898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3565_req_12898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1034), ack => phi_stmt_3565_req_1); -- 
    zeropad3D_cp_element_group_1034: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1034"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1032) & zeropad3D_CP_2152_elements(1033);
      gj_zeropad3D_cp_element_group_1034 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1034), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1035:  transition  input  bypass 
    -- CP-element group 1035: predecessors 
    -- CP-element group 1035: 	500 
    -- CP-element group 1035: successors 
    -- CP-element group 1035: 	1037 
    -- CP-element group 1035:  members (2) 
      -- CP-element group 1035: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3574/SplitProtocol/Sample/$exit
      -- CP-element group 1035: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3574/SplitProtocol/Sample/ra
      -- 
    ra_12915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1035_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3574_inst_ack_0, ack => zeropad3D_CP_2152_elements(1035)); -- 
    -- CP-element group 1036:  transition  input  bypass 
    -- CP-element group 1036: predecessors 
    -- CP-element group 1036: 	500 
    -- CP-element group 1036: successors 
    -- CP-element group 1036: 	1037 
    -- CP-element group 1036:  members (2) 
      -- CP-element group 1036: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3574/SplitProtocol/Update/$exit
      -- CP-element group 1036: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3574/SplitProtocol/Update/ca
      -- 
    ca_12920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1036_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3574_inst_ack_1, ack => zeropad3D_CP_2152_elements(1036)); -- 
    -- CP-element group 1037:  join  transition  output  bypass 
    -- CP-element group 1037: predecessors 
    -- CP-element group 1037: 	1035 
    -- CP-element group 1037: 	1036 
    -- CP-element group 1037: successors 
    -- CP-element group 1037: 	1038 
    -- CP-element group 1037:  members (5) 
      -- CP-element group 1037: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/$exit
      -- CP-element group 1037: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/$exit
      -- CP-element group 1037: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3574/$exit
      -- CP-element group 1037: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3574/SplitProtocol/$exit
      -- CP-element group 1037: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_req
      -- 
    phi_stmt_3571_req_12921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3571_req_12921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1037), ack => phi_stmt_3571_req_0); -- 
    zeropad3D_cp_element_group_1037: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1037"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1035) & zeropad3D_CP_2152_elements(1036);
      gj_zeropad3D_cp_element_group_1037 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1037), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1038:  join  transition  bypass 
    -- CP-element group 1038: predecessors 
    -- CP-element group 1038: 	1031 
    -- CP-element group 1038: 	1034 
    -- CP-element group 1038: 	1037 
    -- CP-element group 1038: successors 
    -- CP-element group 1038: 	1049 
    -- CP-element group 1038:  members (1) 
      -- CP-element group 1038: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1038: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1038"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1031) & zeropad3D_CP_2152_elements(1034) & zeropad3D_CP_2152_elements(1037);
      gj_zeropad3D_cp_element_group_1038 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1038), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1039:  transition  input  bypass 
    -- CP-element group 1039: predecessors 
    -- CP-element group 1039: 	481 
    -- CP-element group 1039: successors 
    -- CP-element group 1039: 	1041 
    -- CP-element group 1039:  members (2) 
      -- CP-element group 1039: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/type_cast_3561/SplitProtocol/Sample/$exit
      -- CP-element group 1039: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/type_cast_3561/SplitProtocol/Sample/ra
      -- 
    ra_12941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1039_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3561_inst_ack_0, ack => zeropad3D_CP_2152_elements(1039)); -- 
    -- CP-element group 1040:  transition  input  bypass 
    -- CP-element group 1040: predecessors 
    -- CP-element group 1040: 	481 
    -- CP-element group 1040: successors 
    -- CP-element group 1040: 	1041 
    -- CP-element group 1040:  members (2) 
      -- CP-element group 1040: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/type_cast_3561/SplitProtocol/Update/$exit
      -- CP-element group 1040: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/type_cast_3561/SplitProtocol/Update/ca
      -- 
    ca_12946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1040_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3561_inst_ack_1, ack => zeropad3D_CP_2152_elements(1040)); -- 
    -- CP-element group 1041:  join  transition  output  bypass 
    -- CP-element group 1041: predecessors 
    -- CP-element group 1041: 	1039 
    -- CP-element group 1041: 	1040 
    -- CP-element group 1041: successors 
    -- CP-element group 1041: 	1048 
    -- CP-element group 1041:  members (5) 
      -- CP-element group 1041: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/$exit
      -- CP-element group 1041: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/$exit
      -- CP-element group 1041: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/type_cast_3561/$exit
      -- CP-element group 1041: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_sources/type_cast_3561/SplitProtocol/$exit
      -- CP-element group 1041: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3558/phi_stmt_3558_req
      -- 
    phi_stmt_3558_req_12947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3558_req_12947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1041), ack => phi_stmt_3558_req_0); -- 
    zeropad3D_cp_element_group_1041: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1041"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1039) & zeropad3D_CP_2152_elements(1040);
      gj_zeropad3D_cp_element_group_1041 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1041), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1042:  transition  input  bypass 
    -- CP-element group 1042: predecessors 
    -- CP-element group 1042: 	481 
    -- CP-element group 1042: successors 
    -- CP-element group 1042: 	1044 
    -- CP-element group 1042:  members (2) 
      -- CP-element group 1042: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3568/SplitProtocol/Sample/$exit
      -- CP-element group 1042: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3568/SplitProtocol/Sample/ra
      -- 
    ra_12964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1042_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3568_inst_ack_0, ack => zeropad3D_CP_2152_elements(1042)); -- 
    -- CP-element group 1043:  transition  input  bypass 
    -- CP-element group 1043: predecessors 
    -- CP-element group 1043: 	481 
    -- CP-element group 1043: successors 
    -- CP-element group 1043: 	1044 
    -- CP-element group 1043:  members (2) 
      -- CP-element group 1043: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3568/SplitProtocol/Update/$exit
      -- CP-element group 1043: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3568/SplitProtocol/Update/ca
      -- 
    ca_12969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1043_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3568_inst_ack_1, ack => zeropad3D_CP_2152_elements(1043)); -- 
    -- CP-element group 1044:  join  transition  output  bypass 
    -- CP-element group 1044: predecessors 
    -- CP-element group 1044: 	1042 
    -- CP-element group 1044: 	1043 
    -- CP-element group 1044: successors 
    -- CP-element group 1044: 	1048 
    -- CP-element group 1044:  members (5) 
      -- CP-element group 1044: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/$exit
      -- CP-element group 1044: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/$exit
      -- CP-element group 1044: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3568/$exit
      -- CP-element group 1044: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_sources/type_cast_3568/SplitProtocol/$exit
      -- CP-element group 1044: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3565/phi_stmt_3565_req
      -- 
    phi_stmt_3565_req_12970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3565_req_12970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1044), ack => phi_stmt_3565_req_0); -- 
    zeropad3D_cp_element_group_1044: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1044"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1042) & zeropad3D_CP_2152_elements(1043);
      gj_zeropad3D_cp_element_group_1044 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1044), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1045:  transition  input  bypass 
    -- CP-element group 1045: predecessors 
    -- CP-element group 1045: 	481 
    -- CP-element group 1045: successors 
    -- CP-element group 1045: 	1047 
    -- CP-element group 1045:  members (2) 
      -- CP-element group 1045: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3576/SplitProtocol/Sample/$exit
      -- CP-element group 1045: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3576/SplitProtocol/Sample/ra
      -- 
    ra_12987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1045_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3576_inst_ack_0, ack => zeropad3D_CP_2152_elements(1045)); -- 
    -- CP-element group 1046:  transition  input  bypass 
    -- CP-element group 1046: predecessors 
    -- CP-element group 1046: 	481 
    -- CP-element group 1046: successors 
    -- CP-element group 1046: 	1047 
    -- CP-element group 1046:  members (2) 
      -- CP-element group 1046: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3576/SplitProtocol/Update/$exit
      -- CP-element group 1046: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3576/SplitProtocol/Update/ca
      -- 
    ca_12992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1046_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3576_inst_ack_1, ack => zeropad3D_CP_2152_elements(1046)); -- 
    -- CP-element group 1047:  join  transition  output  bypass 
    -- CP-element group 1047: predecessors 
    -- CP-element group 1047: 	1045 
    -- CP-element group 1047: 	1046 
    -- CP-element group 1047: successors 
    -- CP-element group 1047: 	1048 
    -- CP-element group 1047:  members (5) 
      -- CP-element group 1047: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/$exit
      -- CP-element group 1047: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/$exit
      -- CP-element group 1047: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3576/$exit
      -- CP-element group 1047: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_sources/type_cast_3576/SplitProtocol/$exit
      -- CP-element group 1047: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3571/phi_stmt_3571_req
      -- 
    phi_stmt_3571_req_12993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3571_req_12993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1047), ack => phi_stmt_3571_req_1); -- 
    zeropad3D_cp_element_group_1047: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1047"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1045) & zeropad3D_CP_2152_elements(1046);
      gj_zeropad3D_cp_element_group_1047 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1047), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1048:  join  transition  bypass 
    -- CP-element group 1048: predecessors 
    -- CP-element group 1048: 	1041 
    -- CP-element group 1048: 	1044 
    -- CP-element group 1048: 	1047 
    -- CP-element group 1048: successors 
    -- CP-element group 1048: 	1049 
    -- CP-element group 1048:  members (1) 
      -- CP-element group 1048: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1048: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1048"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1041) & zeropad3D_CP_2152_elements(1044) & zeropad3D_CP_2152_elements(1047);
      gj_zeropad3D_cp_element_group_1048 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1048), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1049:  merge  fork  transition  place  bypass 
    -- CP-element group 1049: predecessors 
    -- CP-element group 1049: 	1038 
    -- CP-element group 1049: 	1048 
    -- CP-element group 1049: successors 
    -- CP-element group 1049: 	1050 
    -- CP-element group 1049: 	1051 
    -- CP-element group 1049: 	1052 
    -- CP-element group 1049:  members (2) 
      -- CP-element group 1049: 	 branch_block_stmt_714/merge_stmt_3557_PhiReqMerge
      -- CP-element group 1049: 	 branch_block_stmt_714/merge_stmt_3557_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1049) <= OrReduce(zeropad3D_CP_2152_elements(1038) & zeropad3D_CP_2152_elements(1048));
    -- CP-element group 1050:  transition  input  bypass 
    -- CP-element group 1050: predecessors 
    -- CP-element group 1050: 	1049 
    -- CP-element group 1050: successors 
    -- CP-element group 1050: 	1053 
    -- CP-element group 1050:  members (1) 
      -- CP-element group 1050: 	 branch_block_stmt_714/merge_stmt_3557_PhiAck/phi_stmt_3558_ack
      -- 
    phi_stmt_3558_ack_12998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1050_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3558_ack_0, ack => zeropad3D_CP_2152_elements(1050)); -- 
    -- CP-element group 1051:  transition  input  bypass 
    -- CP-element group 1051: predecessors 
    -- CP-element group 1051: 	1049 
    -- CP-element group 1051: successors 
    -- CP-element group 1051: 	1053 
    -- CP-element group 1051:  members (1) 
      -- CP-element group 1051: 	 branch_block_stmt_714/merge_stmt_3557_PhiAck/phi_stmt_3565_ack
      -- 
    phi_stmt_3565_ack_12999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1051_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3565_ack_0, ack => zeropad3D_CP_2152_elements(1051)); -- 
    -- CP-element group 1052:  transition  input  bypass 
    -- CP-element group 1052: predecessors 
    -- CP-element group 1052: 	1049 
    -- CP-element group 1052: successors 
    -- CP-element group 1052: 	1053 
    -- CP-element group 1052:  members (1) 
      -- CP-element group 1052: 	 branch_block_stmt_714/merge_stmt_3557_PhiAck/phi_stmt_3571_ack
      -- 
    phi_stmt_3571_ack_13000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1052_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3571_ack_0, ack => zeropad3D_CP_2152_elements(1052)); -- 
    -- CP-element group 1053:  join  transition  bypass 
    -- CP-element group 1053: predecessors 
    -- CP-element group 1053: 	1050 
    -- CP-element group 1053: 	1051 
    -- CP-element group 1053: 	1052 
    -- CP-element group 1053: successors 
    -- CP-element group 1053: 	5 
    -- CP-element group 1053:  members (1) 
      -- CP-element group 1053: 	 branch_block_stmt_714/merge_stmt_3557_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1053: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1053"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1050) & zeropad3D_CP_2152_elements(1051) & zeropad3D_CP_2152_elements(1052);
      gj_zeropad3D_cp_element_group_1053 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1053), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1054:  transition  input  bypass 
    -- CP-element group 1054: predecessors 
    -- CP-element group 1054: 	499 
    -- CP-element group 1054: successors 
    -- CP-element group 1054: 	1056 
    -- CP-element group 1054:  members (2) 
      -- CP-element group 1054: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/type_cast_3583/SplitProtocol/Sample/$exit
      -- CP-element group 1054: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/type_cast_3583/SplitProtocol/Sample/ra
      -- 
    ra_13020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1054_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3583_inst_ack_0, ack => zeropad3D_CP_2152_elements(1054)); -- 
    -- CP-element group 1055:  transition  input  bypass 
    -- CP-element group 1055: predecessors 
    -- CP-element group 1055: 	499 
    -- CP-element group 1055: successors 
    -- CP-element group 1055: 	1056 
    -- CP-element group 1055:  members (2) 
      -- CP-element group 1055: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/type_cast_3583/SplitProtocol/Update/$exit
      -- CP-element group 1055: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/type_cast_3583/SplitProtocol/Update/ca
      -- 
    ca_13025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1055_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3583_inst_ack_1, ack => zeropad3D_CP_2152_elements(1055)); -- 
    -- CP-element group 1056:  join  transition  output  bypass 
    -- CP-element group 1056: predecessors 
    -- CP-element group 1056: 	1054 
    -- CP-element group 1056: 	1055 
    -- CP-element group 1056: successors 
    -- CP-element group 1056: 	1063 
    -- CP-element group 1056:  members (5) 
      -- CP-element group 1056: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/$exit
      -- CP-element group 1056: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/$exit
      -- CP-element group 1056: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/type_cast_3583/$exit
      -- CP-element group 1056: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_sources/type_cast_3583/SplitProtocol/$exit
      -- CP-element group 1056: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3580/phi_stmt_3580_req
      -- 
    phi_stmt_3580_req_13026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3580_req_13026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1056), ack => phi_stmt_3580_req_0); -- 
    zeropad3D_cp_element_group_1056: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1056"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1054) & zeropad3D_CP_2152_elements(1055);
      gj_zeropad3D_cp_element_group_1056 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1056), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1057:  transition  input  bypass 
    -- CP-element group 1057: predecessors 
    -- CP-element group 1057: 	499 
    -- CP-element group 1057: successors 
    -- CP-element group 1057: 	1059 
    -- CP-element group 1057:  members (2) 
      -- CP-element group 1057: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/type_cast_3587/SplitProtocol/Sample/$exit
      -- CP-element group 1057: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/type_cast_3587/SplitProtocol/Sample/ra
      -- 
    ra_13043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1057_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3587_inst_ack_0, ack => zeropad3D_CP_2152_elements(1057)); -- 
    -- CP-element group 1058:  transition  input  bypass 
    -- CP-element group 1058: predecessors 
    -- CP-element group 1058: 	499 
    -- CP-element group 1058: successors 
    -- CP-element group 1058: 	1059 
    -- CP-element group 1058:  members (2) 
      -- CP-element group 1058: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/type_cast_3587/SplitProtocol/Update/$exit
      -- CP-element group 1058: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/type_cast_3587/SplitProtocol/Update/ca
      -- 
    ca_13048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1058_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3587_inst_ack_1, ack => zeropad3D_CP_2152_elements(1058)); -- 
    -- CP-element group 1059:  join  transition  output  bypass 
    -- CP-element group 1059: predecessors 
    -- CP-element group 1059: 	1057 
    -- CP-element group 1059: 	1058 
    -- CP-element group 1059: successors 
    -- CP-element group 1059: 	1063 
    -- CP-element group 1059:  members (5) 
      -- CP-element group 1059: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/$exit
      -- CP-element group 1059: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/$exit
      -- CP-element group 1059: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/type_cast_3587/$exit
      -- CP-element group 1059: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_sources/type_cast_3587/SplitProtocol/$exit
      -- CP-element group 1059: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3584/phi_stmt_3584_req
      -- 
    phi_stmt_3584_req_13049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3584_req_13049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1059), ack => phi_stmt_3584_req_0); -- 
    zeropad3D_cp_element_group_1059: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1059"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1057) & zeropad3D_CP_2152_elements(1058);
      gj_zeropad3D_cp_element_group_1059 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1059), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1060:  transition  input  bypass 
    -- CP-element group 1060: predecessors 
    -- CP-element group 1060: 	499 
    -- CP-element group 1060: successors 
    -- CP-element group 1060: 	1062 
    -- CP-element group 1060:  members (2) 
      -- CP-element group 1060: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/type_cast_3591/SplitProtocol/Sample/$exit
      -- CP-element group 1060: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/type_cast_3591/SplitProtocol/Sample/ra
      -- 
    ra_13066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1060_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3591_inst_ack_0, ack => zeropad3D_CP_2152_elements(1060)); -- 
    -- CP-element group 1061:  transition  input  bypass 
    -- CP-element group 1061: predecessors 
    -- CP-element group 1061: 	499 
    -- CP-element group 1061: successors 
    -- CP-element group 1061: 	1062 
    -- CP-element group 1061:  members (2) 
      -- CP-element group 1061: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/type_cast_3591/SplitProtocol/Update/$exit
      -- CP-element group 1061: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/type_cast_3591/SplitProtocol/Update/ca
      -- 
    ca_13071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1061_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3591_inst_ack_1, ack => zeropad3D_CP_2152_elements(1061)); -- 
    -- CP-element group 1062:  join  transition  output  bypass 
    -- CP-element group 1062: predecessors 
    -- CP-element group 1062: 	1060 
    -- CP-element group 1062: 	1061 
    -- CP-element group 1062: successors 
    -- CP-element group 1062: 	1063 
    -- CP-element group 1062:  members (5) 
      -- CP-element group 1062: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/$exit
      -- CP-element group 1062: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/$exit
      -- CP-element group 1062: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/type_cast_3591/$exit
      -- CP-element group 1062: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_sources/type_cast_3591/SplitProtocol/$exit
      -- CP-element group 1062: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/phi_stmt_3588/phi_stmt_3588_req
      -- 
    phi_stmt_3588_req_13072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3588_req_13072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1062), ack => phi_stmt_3588_req_0); -- 
    zeropad3D_cp_element_group_1062: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1062"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1060) & zeropad3D_CP_2152_elements(1061);
      gj_zeropad3D_cp_element_group_1062 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1062), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1063:  join  fork  transition  place  bypass 
    -- CP-element group 1063: predecessors 
    -- CP-element group 1063: 	1056 
    -- CP-element group 1063: 	1059 
    -- CP-element group 1063: 	1062 
    -- CP-element group 1063: successors 
    -- CP-element group 1063: 	1064 
    -- CP-element group 1063: 	1065 
    -- CP-element group 1063: 	1066 
    -- CP-element group 1063:  members (3) 
      -- CP-element group 1063: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/$exit
      -- CP-element group 1063: 	 branch_block_stmt_714/merge_stmt_3579_PhiReqMerge
      -- CP-element group 1063: 	 branch_block_stmt_714/merge_stmt_3579_PhiAck/$entry
      -- 
    zeropad3D_cp_element_group_1063: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1063"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1056) & zeropad3D_CP_2152_elements(1059) & zeropad3D_CP_2152_elements(1062);
      gj_zeropad3D_cp_element_group_1063 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1063), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1064:  transition  input  bypass 
    -- CP-element group 1064: predecessors 
    -- CP-element group 1064: 	1063 
    -- CP-element group 1064: successors 
    -- CP-element group 1064: 	1067 
    -- CP-element group 1064:  members (1) 
      -- CP-element group 1064: 	 branch_block_stmt_714/merge_stmt_3579_PhiAck/phi_stmt_3580_ack
      -- 
    phi_stmt_3580_ack_13077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1064_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3580_ack_0, ack => zeropad3D_CP_2152_elements(1064)); -- 
    -- CP-element group 1065:  transition  input  bypass 
    -- CP-element group 1065: predecessors 
    -- CP-element group 1065: 	1063 
    -- CP-element group 1065: successors 
    -- CP-element group 1065: 	1067 
    -- CP-element group 1065:  members (1) 
      -- CP-element group 1065: 	 branch_block_stmt_714/merge_stmt_3579_PhiAck/phi_stmt_3584_ack
      -- 
    phi_stmt_3584_ack_13078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1065_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3584_ack_0, ack => zeropad3D_CP_2152_elements(1065)); -- 
    -- CP-element group 1066:  transition  input  bypass 
    -- CP-element group 1066: predecessors 
    -- CP-element group 1066: 	1063 
    -- CP-element group 1066: successors 
    -- CP-element group 1066: 	1067 
    -- CP-element group 1066:  members (1) 
      -- CP-element group 1066: 	 branch_block_stmt_714/merge_stmt_3579_PhiAck/phi_stmt_3588_ack
      -- 
    phi_stmt_3588_ack_13079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1066_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3588_ack_0, ack => zeropad3D_CP_2152_elements(1066)); -- 
    -- CP-element group 1067:  join  fork  transition  place  output  bypass 
    -- CP-element group 1067: predecessors 
    -- CP-element group 1067: 	1064 
    -- CP-element group 1067: 	1065 
    -- CP-element group 1067: 	1066 
    -- CP-element group 1067: successors 
    -- CP-element group 1067: 	501 
    -- CP-element group 1067: 	502 
    -- CP-element group 1067: 	503 
    -- CP-element group 1067: 	504 
    -- CP-element group 1067: 	505 
    -- CP-element group 1067: 	506 
    -- CP-element group 1067: 	507 
    -- CP-element group 1067: 	508 
    -- CP-element group 1067: 	509 
    -- CP-element group 1067: 	510 
    -- CP-element group 1067: 	511 
    -- CP-element group 1067: 	512 
    -- CP-element group 1067: 	514 
    -- CP-element group 1067: 	516 
    -- CP-element group 1067:  members (98) 
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726__entry__
      -- CP-element group 1067: 	 branch_block_stmt_714/merge_stmt_3579__exit__
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3595_Sample/rr
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3595_Update/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3605_Update/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_update_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3595_Update/cr
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3605_sample_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_sample_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3595_Sample/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3595_update_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3605_Update/cr
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3595_sample_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3605_Sample/rr
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3605_Sample/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3605_update_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_word_address_calculated
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_root_address_calculated
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Sample/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Sample/word_access_start/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Sample/word_access_start/word_0/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Sample/word_access_start/word_0/rr
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Update/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Update/word_access_complete/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Update/word_access_complete/word_0/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_pad_3614_Update/word_access_complete/word_0/cr
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_sample_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_update_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_word_address_calculated
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_root_address_calculated
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Sample/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Sample/word_access_start/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Sample/word_access_start/word_0/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Sample/word_access_start/word_0/rr
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Update/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Update/word_access_complete/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Update/word_access_complete/word_0/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/LOAD_depth_high_3617_Update/word_access_complete/word_0/cr
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_sample_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_update_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_base_address_calculated
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3684_Update/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_word_address_calculated
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_root_address_calculated
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_base_address_resized
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_base_addr_resize/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_base_addr_resize/$exit
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_base_addr_resize/base_resize_req
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_base_addr_resize/base_resize_ack
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_base_plus_offset/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_base_plus_offset/$exit
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_base_plus_offset/sum_rename_req
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_base_plus_offset/sum_rename_ack
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_word_addrgen/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_word_addrgen/$exit
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_word_addrgen/root_register_req
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_word_addrgen/root_register_ack
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Sample/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Sample/word_access_start/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Sample/word_access_start/word_0/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Sample/word_access_start/word_0/rr
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Update/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Update/word_access_complete/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Update/word_access_complete/word_0/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3629_Update/word_access_complete/word_0/cr
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_sample_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_update_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_base_address_calculated
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_word_address_calculated
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_root_address_calculated
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_base_address_resized
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_base_addr_resize/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_base_addr_resize/$exit
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_base_addr_resize/base_resize_req
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_base_addr_resize/base_resize_ack
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_base_plus_offset/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_base_plus_offset/$exit
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_base_plus_offset/sum_rename_req
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_base_plus_offset/sum_rename_ack
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_word_addrgen/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_word_addrgen/$exit
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_word_addrgen/root_register_req
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_word_addrgen/root_register_ack
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Sample/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Sample/word_access_start/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Sample/word_access_start/word_0/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Sample/word_access_start/word_0/rr
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Update/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Update/word_access_complete/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Update/word_access_complete/word_0/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/ptr_deref_3641_Update/word_access_complete/word_0/cr
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3645_update_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3645_Update/$entry
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3645_Update/cr
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3684_update_start_
      -- CP-element group 1067: 	 branch_block_stmt_714/assign_stmt_3596_to_assign_stmt_3726/type_cast_3684_Update/cr
      -- CP-element group 1067: 	 branch_block_stmt_714/merge_stmt_3579_PhiAck/$exit
      -- 
    rr_7949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => type_cast_3595_inst_req_0); -- 
    cr_7954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => type_cast_3595_inst_req_1); -- 
    cr_7968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => type_cast_3605_inst_req_1); -- 
    rr_7963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => type_cast_3605_inst_req_0); -- 
    rr_7985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => LOAD_pad_3614_load_0_req_0); -- 
    cr_7996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => LOAD_pad_3614_load_0_req_1); -- 
    rr_8018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => LOAD_depth_high_3617_load_0_req_0); -- 
    cr_8029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => LOAD_depth_high_3617_load_0_req_1); -- 
    rr_8068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => ptr_deref_3629_load_0_req_0); -- 
    cr_8079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => ptr_deref_3629_load_0_req_1); -- 
    rr_8118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => ptr_deref_3641_load_0_req_0); -- 
    cr_8129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => ptr_deref_3641_load_0_req_1); -- 
    cr_8148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => type_cast_3645_inst_req_1); -- 
    cr_8162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1067), ack => type_cast_3684_inst_req_1); -- 
    zeropad3D_cp_element_group_1067: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1067"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1064) & zeropad3D_CP_2152_elements(1065) & zeropad3D_CP_2152_elements(1066);
      gj_zeropad3D_cp_element_group_1067 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1067), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1068:  transition  input  bypass 
    -- CP-element group 1068: predecessors 
    -- CP-element group 1068: 	6 
    -- CP-element group 1068: successors 
    -- CP-element group 1068: 	1070 
    -- CP-element group 1068:  members (2) 
      -- CP-element group 1068: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/type_cast_3732/SplitProtocol/Sample/$exit
      -- CP-element group 1068: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/type_cast_3732/SplitProtocol/Sample/ra
      -- 
    ra_13099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1068_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3732_inst_ack_0, ack => zeropad3D_CP_2152_elements(1068)); -- 
    -- CP-element group 1069:  transition  input  bypass 
    -- CP-element group 1069: predecessors 
    -- CP-element group 1069: 	6 
    -- CP-element group 1069: successors 
    -- CP-element group 1069: 	1070 
    -- CP-element group 1069:  members (2) 
      -- CP-element group 1069: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/type_cast_3732/SplitProtocol/Update/$exit
      -- CP-element group 1069: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/type_cast_3732/SplitProtocol/Update/ca
      -- 
    ca_13104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1069_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3732_inst_ack_1, ack => zeropad3D_CP_2152_elements(1069)); -- 
    -- CP-element group 1070:  join  transition  output  bypass 
    -- CP-element group 1070: predecessors 
    -- CP-element group 1070: 	1068 
    -- CP-element group 1070: 	1069 
    -- CP-element group 1070: successors 
    -- CP-element group 1070: 	1077 
    -- CP-element group 1070:  members (5) 
      -- CP-element group 1070: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/$exit
      -- CP-element group 1070: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/$exit
      -- CP-element group 1070: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/type_cast_3732/$exit
      -- CP-element group 1070: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/type_cast_3732/SplitProtocol/$exit
      -- CP-element group 1070: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_req
      -- 
    phi_stmt_3729_req_13105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3729_req_13105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1070), ack => phi_stmt_3729_req_0); -- 
    zeropad3D_cp_element_group_1070: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1070"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1068) & zeropad3D_CP_2152_elements(1069);
      gj_zeropad3D_cp_element_group_1070 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1070), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1071:  transition  input  bypass 
    -- CP-element group 1071: predecessors 
    -- CP-element group 1071: 	6 
    -- CP-element group 1071: successors 
    -- CP-element group 1071: 	1073 
    -- CP-element group 1071:  members (2) 
      -- CP-element group 1071: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3739/SplitProtocol/Sample/$exit
      -- CP-element group 1071: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3739/SplitProtocol/Sample/ra
      -- 
    ra_13122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1071_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3739_inst_ack_0, ack => zeropad3D_CP_2152_elements(1071)); -- 
    -- CP-element group 1072:  transition  input  bypass 
    -- CP-element group 1072: predecessors 
    -- CP-element group 1072: 	6 
    -- CP-element group 1072: successors 
    -- CP-element group 1072: 	1073 
    -- CP-element group 1072:  members (2) 
      -- CP-element group 1072: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3739/SplitProtocol/Update/$exit
      -- CP-element group 1072: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3739/SplitProtocol/Update/ca
      -- 
    ca_13127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1072_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3739_inst_ack_1, ack => zeropad3D_CP_2152_elements(1072)); -- 
    -- CP-element group 1073:  join  transition  output  bypass 
    -- CP-element group 1073: predecessors 
    -- CP-element group 1073: 	1071 
    -- CP-element group 1073: 	1072 
    -- CP-element group 1073: successors 
    -- CP-element group 1073: 	1077 
    -- CP-element group 1073:  members (5) 
      -- CP-element group 1073: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/$exit
      -- CP-element group 1073: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/$exit
      -- CP-element group 1073: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3739/$exit
      -- CP-element group 1073: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3739/SplitProtocol/$exit
      -- CP-element group 1073: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_req
      -- 
    phi_stmt_3736_req_13128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3736_req_13128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1073), ack => phi_stmt_3736_req_0); -- 
    zeropad3D_cp_element_group_1073: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1073"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1071) & zeropad3D_CP_2152_elements(1072);
      gj_zeropad3D_cp_element_group_1073 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1073), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1074:  transition  input  bypass 
    -- CP-element group 1074: predecessors 
    -- CP-element group 1074: 	6 
    -- CP-element group 1074: successors 
    -- CP-element group 1074: 	1076 
    -- CP-element group 1074:  members (2) 
      -- CP-element group 1074: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3747/SplitProtocol/Sample/$exit
      -- CP-element group 1074: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3747/SplitProtocol/Sample/ra
      -- 
    ra_13145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1074_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3747_inst_ack_0, ack => zeropad3D_CP_2152_elements(1074)); -- 
    -- CP-element group 1075:  transition  input  bypass 
    -- CP-element group 1075: predecessors 
    -- CP-element group 1075: 	6 
    -- CP-element group 1075: successors 
    -- CP-element group 1075: 	1076 
    -- CP-element group 1075:  members (2) 
      -- CP-element group 1075: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3747/SplitProtocol/Update/$exit
      -- CP-element group 1075: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3747/SplitProtocol/Update/ca
      -- 
    ca_13150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1075_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3747_inst_ack_1, ack => zeropad3D_CP_2152_elements(1075)); -- 
    -- CP-element group 1076:  join  transition  output  bypass 
    -- CP-element group 1076: predecessors 
    -- CP-element group 1076: 	1074 
    -- CP-element group 1076: 	1075 
    -- CP-element group 1076: successors 
    -- CP-element group 1076: 	1077 
    -- CP-element group 1076:  members (5) 
      -- CP-element group 1076: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/$exit
      -- CP-element group 1076: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/$exit
      -- CP-element group 1076: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3747/$exit
      -- CP-element group 1076: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3747/SplitProtocol/$exit
      -- CP-element group 1076: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_req
      -- 
    phi_stmt_3742_req_13151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3742_req_13151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1076), ack => phi_stmt_3742_req_1); -- 
    zeropad3D_cp_element_group_1076: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1076"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1074) & zeropad3D_CP_2152_elements(1075);
      gj_zeropad3D_cp_element_group_1076 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1076), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1077:  join  transition  bypass 
    -- CP-element group 1077: predecessors 
    -- CP-element group 1077: 	1070 
    -- CP-element group 1077: 	1073 
    -- CP-element group 1077: 	1076 
    -- CP-element group 1077: successors 
    -- CP-element group 1077: 	1086 
    -- CP-element group 1077:  members (1) 
      -- CP-element group 1077: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1077: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1077"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1070) & zeropad3D_CP_2152_elements(1073) & zeropad3D_CP_2152_elements(1076);
      gj_zeropad3D_cp_element_group_1077 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1077), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1078:  transition  output  delay-element  bypass 
    -- CP-element group 1078: predecessors 
    -- CP-element group 1078: 	517 
    -- CP-element group 1078: successors 
    -- CP-element group 1078: 	1085 
    -- CP-element group 1078:  members (4) 
      -- CP-element group 1078: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3729/$exit
      -- CP-element group 1078: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/$exit
      -- CP-element group 1078: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_sources/type_cast_3735_konst_delay_trans
      -- CP-element group 1078: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3729/phi_stmt_3729_req
      -- 
    phi_stmt_3729_req_13162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3729_req_13162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1078), ack => phi_stmt_3729_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(1078) is a control-delay.
    cp_element_1078_delay: control_delay_element  generic map(name => " 1078_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(517), ack => zeropad3D_CP_2152_elements(1078), clk => clk, reset =>reset);
    -- CP-element group 1079:  transition  input  bypass 
    -- CP-element group 1079: predecessors 
    -- CP-element group 1079: 	517 
    -- CP-element group 1079: successors 
    -- CP-element group 1079: 	1081 
    -- CP-element group 1079:  members (2) 
      -- CP-element group 1079: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3741/SplitProtocol/Sample/$exit
      -- CP-element group 1079: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3741/SplitProtocol/Sample/ra
      -- 
    ra_13179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1079_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3741_inst_ack_0, ack => zeropad3D_CP_2152_elements(1079)); -- 
    -- CP-element group 1080:  transition  input  bypass 
    -- CP-element group 1080: predecessors 
    -- CP-element group 1080: 	517 
    -- CP-element group 1080: successors 
    -- CP-element group 1080: 	1081 
    -- CP-element group 1080:  members (2) 
      -- CP-element group 1080: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3741/SplitProtocol/Update/$exit
      -- CP-element group 1080: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3741/SplitProtocol/Update/ca
      -- 
    ca_13184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1080_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3741_inst_ack_1, ack => zeropad3D_CP_2152_elements(1080)); -- 
    -- CP-element group 1081:  join  transition  output  bypass 
    -- CP-element group 1081: predecessors 
    -- CP-element group 1081: 	1079 
    -- CP-element group 1081: 	1080 
    -- CP-element group 1081: successors 
    -- CP-element group 1081: 	1085 
    -- CP-element group 1081:  members (5) 
      -- CP-element group 1081: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/$exit
      -- CP-element group 1081: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/$exit
      -- CP-element group 1081: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3741/$exit
      -- CP-element group 1081: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_sources/type_cast_3741/SplitProtocol/$exit
      -- CP-element group 1081: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3736/phi_stmt_3736_req
      -- 
    phi_stmt_3736_req_13185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3736_req_13185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1081), ack => phi_stmt_3736_req_1); -- 
    zeropad3D_cp_element_group_1081: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1081"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1079) & zeropad3D_CP_2152_elements(1080);
      gj_zeropad3D_cp_element_group_1081 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1081), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1082:  transition  input  bypass 
    -- CP-element group 1082: predecessors 
    -- CP-element group 1082: 	517 
    -- CP-element group 1082: successors 
    -- CP-element group 1082: 	1084 
    -- CP-element group 1082:  members (2) 
      -- CP-element group 1082: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3745/SplitProtocol/Sample/$exit
      -- CP-element group 1082: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3745/SplitProtocol/Sample/ra
      -- 
    ra_13202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1082_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3745_inst_ack_0, ack => zeropad3D_CP_2152_elements(1082)); -- 
    -- CP-element group 1083:  transition  input  bypass 
    -- CP-element group 1083: predecessors 
    -- CP-element group 1083: 	517 
    -- CP-element group 1083: successors 
    -- CP-element group 1083: 	1084 
    -- CP-element group 1083:  members (2) 
      -- CP-element group 1083: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3745/SplitProtocol/Update/$exit
      -- CP-element group 1083: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3745/SplitProtocol/Update/ca
      -- 
    ca_13207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1083_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3745_inst_ack_1, ack => zeropad3D_CP_2152_elements(1083)); -- 
    -- CP-element group 1084:  join  transition  output  bypass 
    -- CP-element group 1084: predecessors 
    -- CP-element group 1084: 	1082 
    -- CP-element group 1084: 	1083 
    -- CP-element group 1084: successors 
    -- CP-element group 1084: 	1085 
    -- CP-element group 1084:  members (5) 
      -- CP-element group 1084: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/$exit
      -- CP-element group 1084: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/$exit
      -- CP-element group 1084: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3745/$exit
      -- CP-element group 1084: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_sources/type_cast_3745/SplitProtocol/$exit
      -- CP-element group 1084: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3742/phi_stmt_3742_req
      -- 
    phi_stmt_3742_req_13208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3742_req_13208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1084), ack => phi_stmt_3742_req_0); -- 
    zeropad3D_cp_element_group_1084: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1084"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1082) & zeropad3D_CP_2152_elements(1083);
      gj_zeropad3D_cp_element_group_1084 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1084), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1085:  join  transition  bypass 
    -- CP-element group 1085: predecessors 
    -- CP-element group 1085: 	1078 
    -- CP-element group 1085: 	1081 
    -- CP-element group 1085: 	1084 
    -- CP-element group 1085: successors 
    -- CP-element group 1085: 	1086 
    -- CP-element group 1085:  members (1) 
      -- CP-element group 1085: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1085: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1085"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1078) & zeropad3D_CP_2152_elements(1081) & zeropad3D_CP_2152_elements(1084);
      gj_zeropad3D_cp_element_group_1085 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1085), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1086:  merge  fork  transition  place  bypass 
    -- CP-element group 1086: predecessors 
    -- CP-element group 1086: 	1077 
    -- CP-element group 1086: 	1085 
    -- CP-element group 1086: successors 
    -- CP-element group 1086: 	1087 
    -- CP-element group 1086: 	1088 
    -- CP-element group 1086: 	1089 
    -- CP-element group 1086:  members (2) 
      -- CP-element group 1086: 	 branch_block_stmt_714/merge_stmt_3728_PhiReqMerge
      -- CP-element group 1086: 	 branch_block_stmt_714/merge_stmt_3728_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1086) <= OrReduce(zeropad3D_CP_2152_elements(1077) & zeropad3D_CP_2152_elements(1085));
    -- CP-element group 1087:  transition  input  bypass 
    -- CP-element group 1087: predecessors 
    -- CP-element group 1087: 	1086 
    -- CP-element group 1087: successors 
    -- CP-element group 1087: 	1090 
    -- CP-element group 1087:  members (1) 
      -- CP-element group 1087: 	 branch_block_stmt_714/merge_stmt_3728_PhiAck/phi_stmt_3729_ack
      -- 
    phi_stmt_3729_ack_13213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1087_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3729_ack_0, ack => zeropad3D_CP_2152_elements(1087)); -- 
    -- CP-element group 1088:  transition  input  bypass 
    -- CP-element group 1088: predecessors 
    -- CP-element group 1088: 	1086 
    -- CP-element group 1088: successors 
    -- CP-element group 1088: 	1090 
    -- CP-element group 1088:  members (1) 
      -- CP-element group 1088: 	 branch_block_stmt_714/merge_stmt_3728_PhiAck/phi_stmt_3736_ack
      -- 
    phi_stmt_3736_ack_13214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1088_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3736_ack_0, ack => zeropad3D_CP_2152_elements(1088)); -- 
    -- CP-element group 1089:  transition  input  bypass 
    -- CP-element group 1089: predecessors 
    -- CP-element group 1089: 	1086 
    -- CP-element group 1089: successors 
    -- CP-element group 1089: 	1090 
    -- CP-element group 1089:  members (1) 
      -- CP-element group 1089: 	 branch_block_stmt_714/merge_stmt_3728_PhiAck/phi_stmt_3742_ack
      -- 
    phi_stmt_3742_ack_13215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1089_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3742_ack_0, ack => zeropad3D_CP_2152_elements(1089)); -- 
    -- CP-element group 1090:  join  fork  transition  place  output  bypass 
    -- CP-element group 1090: predecessors 
    -- CP-element group 1090: 	1087 
    -- CP-element group 1090: 	1088 
    -- CP-element group 1090: 	1089 
    -- CP-element group 1090: successors 
    -- CP-element group 1090: 	518 
    -- CP-element group 1090: 	519 
    -- CP-element group 1090:  members (10) 
      -- CP-element group 1090: 	 branch_block_stmt_714/merge_stmt_3728__exit__
      -- CP-element group 1090: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760__entry__
      -- CP-element group 1090: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/$entry
      -- CP-element group 1090: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/type_cast_3752_sample_start_
      -- CP-element group 1090: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/type_cast_3752_update_start_
      -- CP-element group 1090: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/type_cast_3752_Sample/$entry
      -- CP-element group 1090: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/type_cast_3752_Sample/rr
      -- CP-element group 1090: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/type_cast_3752_Update/$entry
      -- CP-element group 1090: 	 branch_block_stmt_714/assign_stmt_3753_to_assign_stmt_3760/type_cast_3752_Update/cr
      -- CP-element group 1090: 	 branch_block_stmt_714/merge_stmt_3728_PhiAck/$exit
      -- 
    rr_8174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1090), ack => type_cast_3752_inst_req_0); -- 
    cr_8179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1090), ack => type_cast_3752_inst_req_1); -- 
    zeropad3D_cp_element_group_1090: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1090"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1087) & zeropad3D_CP_2152_elements(1088) & zeropad3D_CP_2152_elements(1089);
      gj_zeropad3D_cp_element_group_1090 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1090), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1091:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1091: predecessors 
    -- CP-element group 1091: 	520 
    -- CP-element group 1091: 	527 
    -- CP-element group 1091: 	530 
    -- CP-element group 1091: 	537 
    -- CP-element group 1091: successors 
    -- CP-element group 1091: 	538 
    -- CP-element group 1091: 	539 
    -- CP-element group 1091: 	540 
    -- CP-element group 1091: 	541 
    -- CP-element group 1091: 	544 
    -- CP-element group 1091: 	546 
    -- CP-element group 1091: 	548 
    -- CP-element group 1091: 	550 
    -- CP-element group 1091:  members (33) 
      -- CP-element group 1091: 	 branch_block_stmt_714/merge_stmt_3850__exit__
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906__entry__
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/$entry
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3854_sample_start_
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3854_update_start_
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3854_Sample/$entry
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3854_Sample/rr
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3854_Update/$entry
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3854_Update/cr
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3859_sample_start_
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3859_update_start_
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3859_Sample/$entry
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3859_Sample/rr
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3859_Update/$entry
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3859_Update/cr
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3893_update_start_
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3893_Update/$entry
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/type_cast_3893_Update/cr
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/addr_of_3900_update_start_
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_final_index_sum_regn_update_start
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_final_index_sum_regn_Update/$entry
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/array_obj_ref_3899_final_index_sum_regn_Update/req
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/addr_of_3900_complete/$entry
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/addr_of_3900_complete/req
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_update_start_
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Update/$entry
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Update/word_access_complete/$entry
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Update/word_access_complete/word_0/$entry
      -- CP-element group 1091: 	 branch_block_stmt_714/assign_stmt_3855_to_assign_stmt_3906/ptr_deref_3903_Update/word_access_complete/word_0/cr
      -- CP-element group 1091: 	 branch_block_stmt_714/merge_stmt_3850_PhiReqMerge
      -- CP-element group 1091: 	 branch_block_stmt_714/merge_stmt_3850_PhiAck/$entry
      -- CP-element group 1091: 	 branch_block_stmt_714/merge_stmt_3850_PhiAck/$exit
      -- CP-element group 1091: 	 branch_block_stmt_714/merge_stmt_3850_PhiAck/dummy
      -- 
    rr_8384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1091), ack => type_cast_3854_inst_req_0); -- 
    cr_8389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1091), ack => type_cast_3854_inst_req_1); -- 
    rr_8398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1091), ack => type_cast_3859_inst_req_0); -- 
    cr_8403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1091), ack => type_cast_3859_inst_req_1); -- 
    cr_8417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1091), ack => type_cast_3893_inst_req_1); -- 
    req_8448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1091), ack => array_obj_ref_3899_index_offset_req_1); -- 
    req_8463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1091), ack => addr_of_3900_final_reg_req_1); -- 
    cr_8513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1091), ack => ptr_deref_3903_store_0_req_1); -- 
    zeropad3D_CP_2152_elements(1091) <= OrReduce(zeropad3D_CP_2152_elements(520) & zeropad3D_CP_2152_elements(527) & zeropad3D_CP_2152_elements(530) & zeropad3D_CP_2152_elements(537));
    -- CP-element group 1092:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1092: predecessors 
    -- CP-element group 1092: 	551 
    -- CP-element group 1092: 	571 
    -- CP-element group 1092: successors 
    -- CP-element group 1092: 	572 
    -- CP-element group 1092: 	573 
    -- CP-element group 1092:  members (13) 
      -- CP-element group 1092: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033__entry__
      -- CP-element group 1092: 	 branch_block_stmt_714/merge_stmt_4015__exit__
      -- CP-element group 1092: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/type_cast_4019_Update/$entry
      -- CP-element group 1092: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/type_cast_4019_Update/cr
      -- CP-element group 1092: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/type_cast_4019_Sample/rr
      -- CP-element group 1092: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/type_cast_4019_Sample/$entry
      -- CP-element group 1092: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/type_cast_4019_update_start_
      -- CP-element group 1092: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/type_cast_4019_sample_start_
      -- CP-element group 1092: 	 branch_block_stmt_714/assign_stmt_4020_to_assign_stmt_4033/$entry
      -- CP-element group 1092: 	 branch_block_stmt_714/merge_stmt_4015_PhiReqMerge
      -- CP-element group 1092: 	 branch_block_stmt_714/merge_stmt_4015_PhiAck/$entry
      -- CP-element group 1092: 	 branch_block_stmt_714/merge_stmt_4015_PhiAck/$exit
      -- CP-element group 1092: 	 branch_block_stmt_714/merge_stmt_4015_PhiAck/dummy
      -- 
    cr_8767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1092), ack => type_cast_4019_inst_req_1); -- 
    rr_8762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1092), ack => type_cast_4019_inst_req_0); -- 
    zeropad3D_CP_2152_elements(1092) <= OrReduce(zeropad3D_CP_2152_elements(551) & zeropad3D_CP_2152_elements(571));
    -- CP-element group 1093:  transition  output  delay-element  bypass 
    -- CP-element group 1093: predecessors 
    -- CP-element group 1093: 	593 
    -- CP-element group 1093: successors 
    -- CP-element group 1093: 	1100 
    -- CP-element group 1093:  members (4) 
      -- CP-element group 1093: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4133/$exit
      -- CP-element group 1093: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/$exit
      -- CP-element group 1093: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/type_cast_4139_konst_delay_trans
      -- CP-element group 1093: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_req
      -- 
    phi_stmt_4133_req_13326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4133_req_13326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1093), ack => phi_stmt_4133_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(1093) is a control-delay.
    cp_element_1093_delay: control_delay_element  generic map(name => " 1093_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(593), ack => zeropad3D_CP_2152_elements(1093), clk => clk, reset =>reset);
    -- CP-element group 1094:  transition  input  bypass 
    -- CP-element group 1094: predecessors 
    -- CP-element group 1094: 	593 
    -- CP-element group 1094: successors 
    -- CP-element group 1094: 	1096 
    -- CP-element group 1094:  members (2) 
      -- CP-element group 1094: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4145/SplitProtocol/Sample/$exit
      -- CP-element group 1094: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4145/SplitProtocol/Sample/ra
      -- 
    ra_13343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1094_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4145_inst_ack_0, ack => zeropad3D_CP_2152_elements(1094)); -- 
    -- CP-element group 1095:  transition  input  bypass 
    -- CP-element group 1095: predecessors 
    -- CP-element group 1095: 	593 
    -- CP-element group 1095: successors 
    -- CP-element group 1095: 	1096 
    -- CP-element group 1095:  members (2) 
      -- CP-element group 1095: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4145/SplitProtocol/Update/$exit
      -- CP-element group 1095: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4145/SplitProtocol/Update/ca
      -- 
    ca_13348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1095_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4145_inst_ack_1, ack => zeropad3D_CP_2152_elements(1095)); -- 
    -- CP-element group 1096:  join  transition  output  bypass 
    -- CP-element group 1096: predecessors 
    -- CP-element group 1096: 	1094 
    -- CP-element group 1096: 	1095 
    -- CP-element group 1096: successors 
    -- CP-element group 1096: 	1100 
    -- CP-element group 1096:  members (5) 
      -- CP-element group 1096: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/$exit
      -- CP-element group 1096: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/$exit
      -- CP-element group 1096: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4145/$exit
      -- CP-element group 1096: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4145/SplitProtocol/$exit
      -- CP-element group 1096: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_req
      -- 
    phi_stmt_4140_req_13349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4140_req_13349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1096), ack => phi_stmt_4140_req_1); -- 
    zeropad3D_cp_element_group_1096: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1096"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1094) & zeropad3D_CP_2152_elements(1095);
      gj_zeropad3D_cp_element_group_1096 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1096), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1097:  transition  input  bypass 
    -- CP-element group 1097: predecessors 
    -- CP-element group 1097: 	593 
    -- CP-element group 1097: successors 
    -- CP-element group 1097: 	1099 
    -- CP-element group 1097:  members (2) 
      -- CP-element group 1097: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4151/SplitProtocol/Sample/$exit
      -- CP-element group 1097: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4151/SplitProtocol/Sample/ra
      -- 
    ra_13366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1097_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4151_inst_ack_0, ack => zeropad3D_CP_2152_elements(1097)); -- 
    -- CP-element group 1098:  transition  input  bypass 
    -- CP-element group 1098: predecessors 
    -- CP-element group 1098: 	593 
    -- CP-element group 1098: successors 
    -- CP-element group 1098: 	1099 
    -- CP-element group 1098:  members (2) 
      -- CP-element group 1098: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4151/SplitProtocol/Update/$exit
      -- CP-element group 1098: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4151/SplitProtocol/Update/ca
      -- 
    ca_13371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1098_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4151_inst_ack_1, ack => zeropad3D_CP_2152_elements(1098)); -- 
    -- CP-element group 1099:  join  transition  output  bypass 
    -- CP-element group 1099: predecessors 
    -- CP-element group 1099: 	1097 
    -- CP-element group 1099: 	1098 
    -- CP-element group 1099: successors 
    -- CP-element group 1099: 	1100 
    -- CP-element group 1099:  members (5) 
      -- CP-element group 1099: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/$exit
      -- CP-element group 1099: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/$exit
      -- CP-element group 1099: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4151/$exit
      -- CP-element group 1099: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4151/SplitProtocol/$exit
      -- CP-element group 1099: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_req
      -- 
    phi_stmt_4146_req_13372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4146_req_13372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1099), ack => phi_stmt_4146_req_1); -- 
    zeropad3D_cp_element_group_1099: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1099"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1097) & zeropad3D_CP_2152_elements(1098);
      gj_zeropad3D_cp_element_group_1099 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1099), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1100:  join  transition  bypass 
    -- CP-element group 1100: predecessors 
    -- CP-element group 1100: 	1093 
    -- CP-element group 1100: 	1096 
    -- CP-element group 1100: 	1099 
    -- CP-element group 1100: successors 
    -- CP-element group 1100: 	1111 
    -- CP-element group 1100:  members (1) 
      -- CP-element group 1100: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1100: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1100"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1093) & zeropad3D_CP_2152_elements(1096) & zeropad3D_CP_2152_elements(1099);
      gj_zeropad3D_cp_element_group_1100 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1101:  transition  input  bypass 
    -- CP-element group 1101: predecessors 
    -- CP-element group 1101: 	574 
    -- CP-element group 1101: successors 
    -- CP-element group 1101: 	1103 
    -- CP-element group 1101:  members (2) 
      -- CP-element group 1101: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/type_cast_4136/SplitProtocol/Sample/$exit
      -- CP-element group 1101: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/type_cast_4136/SplitProtocol/Sample/ra
      -- 
    ra_13392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4136_inst_ack_0, ack => zeropad3D_CP_2152_elements(1101)); -- 
    -- CP-element group 1102:  transition  input  bypass 
    -- CP-element group 1102: predecessors 
    -- CP-element group 1102: 	574 
    -- CP-element group 1102: successors 
    -- CP-element group 1102: 	1103 
    -- CP-element group 1102:  members (2) 
      -- CP-element group 1102: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/type_cast_4136/SplitProtocol/Update/$exit
      -- CP-element group 1102: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/type_cast_4136/SplitProtocol/Update/ca
      -- 
    ca_13397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4136_inst_ack_1, ack => zeropad3D_CP_2152_elements(1102)); -- 
    -- CP-element group 1103:  join  transition  output  bypass 
    -- CP-element group 1103: predecessors 
    -- CP-element group 1103: 	1101 
    -- CP-element group 1103: 	1102 
    -- CP-element group 1103: successors 
    -- CP-element group 1103: 	1110 
    -- CP-element group 1103:  members (5) 
      -- CP-element group 1103: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/$exit
      -- CP-element group 1103: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/$exit
      -- CP-element group 1103: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/type_cast_4136/$exit
      -- CP-element group 1103: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_sources/type_cast_4136/SplitProtocol/$exit
      -- CP-element group 1103: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4133/phi_stmt_4133_req
      -- 
    phi_stmt_4133_req_13398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4133_req_13398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1103), ack => phi_stmt_4133_req_0); -- 
    zeropad3D_cp_element_group_1103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1101) & zeropad3D_CP_2152_elements(1102);
      gj_zeropad3D_cp_element_group_1103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1104:  transition  input  bypass 
    -- CP-element group 1104: predecessors 
    -- CP-element group 1104: 	574 
    -- CP-element group 1104: successors 
    -- CP-element group 1104: 	1106 
    -- CP-element group 1104:  members (2) 
      -- CP-element group 1104: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4143/SplitProtocol/Sample/$exit
      -- CP-element group 1104: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4143/SplitProtocol/Sample/ra
      -- 
    ra_13415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4143_inst_ack_0, ack => zeropad3D_CP_2152_elements(1104)); -- 
    -- CP-element group 1105:  transition  input  bypass 
    -- CP-element group 1105: predecessors 
    -- CP-element group 1105: 	574 
    -- CP-element group 1105: successors 
    -- CP-element group 1105: 	1106 
    -- CP-element group 1105:  members (2) 
      -- CP-element group 1105: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4143/SplitProtocol/Update/$exit
      -- CP-element group 1105: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4143/SplitProtocol/Update/ca
      -- 
    ca_13420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4143_inst_ack_1, ack => zeropad3D_CP_2152_elements(1105)); -- 
    -- CP-element group 1106:  join  transition  output  bypass 
    -- CP-element group 1106: predecessors 
    -- CP-element group 1106: 	1104 
    -- CP-element group 1106: 	1105 
    -- CP-element group 1106: successors 
    -- CP-element group 1106: 	1110 
    -- CP-element group 1106:  members (5) 
      -- CP-element group 1106: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/$exit
      -- CP-element group 1106: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/$exit
      -- CP-element group 1106: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4143/$exit
      -- CP-element group 1106: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_sources/type_cast_4143/SplitProtocol/$exit
      -- CP-element group 1106: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4140/phi_stmt_4140_req
      -- 
    phi_stmt_4140_req_13421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4140_req_13421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1106), ack => phi_stmt_4140_req_0); -- 
    zeropad3D_cp_element_group_1106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1104) & zeropad3D_CP_2152_elements(1105);
      gj_zeropad3D_cp_element_group_1106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1107:  transition  input  bypass 
    -- CP-element group 1107: predecessors 
    -- CP-element group 1107: 	574 
    -- CP-element group 1107: successors 
    -- CP-element group 1107: 	1109 
    -- CP-element group 1107:  members (2) 
      -- CP-element group 1107: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4149/SplitProtocol/Sample/$exit
      -- CP-element group 1107: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4149/SplitProtocol/Sample/ra
      -- 
    ra_13438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4149_inst_ack_0, ack => zeropad3D_CP_2152_elements(1107)); -- 
    -- CP-element group 1108:  transition  input  bypass 
    -- CP-element group 1108: predecessors 
    -- CP-element group 1108: 	574 
    -- CP-element group 1108: successors 
    -- CP-element group 1108: 	1109 
    -- CP-element group 1108:  members (2) 
      -- CP-element group 1108: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4149/SplitProtocol/Update/$exit
      -- CP-element group 1108: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4149/SplitProtocol/Update/ca
      -- 
    ca_13443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4149_inst_ack_1, ack => zeropad3D_CP_2152_elements(1108)); -- 
    -- CP-element group 1109:  join  transition  output  bypass 
    -- CP-element group 1109: predecessors 
    -- CP-element group 1109: 	1107 
    -- CP-element group 1109: 	1108 
    -- CP-element group 1109: successors 
    -- CP-element group 1109: 	1110 
    -- CP-element group 1109:  members (5) 
      -- CP-element group 1109: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/$exit
      -- CP-element group 1109: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/$exit
      -- CP-element group 1109: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4149/$exit
      -- CP-element group 1109: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_sources/type_cast_4149/SplitProtocol/$exit
      -- CP-element group 1109: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4146/phi_stmt_4146_req
      -- 
    phi_stmt_4146_req_13444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4146_req_13444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1109), ack => phi_stmt_4146_req_0); -- 
    zeropad3D_cp_element_group_1109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1107) & zeropad3D_CP_2152_elements(1108);
      gj_zeropad3D_cp_element_group_1109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1110:  join  transition  bypass 
    -- CP-element group 1110: predecessors 
    -- CP-element group 1110: 	1103 
    -- CP-element group 1110: 	1106 
    -- CP-element group 1110: 	1109 
    -- CP-element group 1110: successors 
    -- CP-element group 1110: 	1111 
    -- CP-element group 1110:  members (1) 
      -- CP-element group 1110: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1103) & zeropad3D_CP_2152_elements(1106) & zeropad3D_CP_2152_elements(1109);
      gj_zeropad3D_cp_element_group_1110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1111:  merge  fork  transition  place  bypass 
    -- CP-element group 1111: predecessors 
    -- CP-element group 1111: 	1100 
    -- CP-element group 1111: 	1110 
    -- CP-element group 1111: successors 
    -- CP-element group 1111: 	1112 
    -- CP-element group 1111: 	1113 
    -- CP-element group 1111: 	1114 
    -- CP-element group 1111:  members (2) 
      -- CP-element group 1111: 	 branch_block_stmt_714/merge_stmt_4132_PhiReqMerge
      -- CP-element group 1111: 	 branch_block_stmt_714/merge_stmt_4132_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1111) <= OrReduce(zeropad3D_CP_2152_elements(1100) & zeropad3D_CP_2152_elements(1110));
    -- CP-element group 1112:  transition  input  bypass 
    -- CP-element group 1112: predecessors 
    -- CP-element group 1112: 	1111 
    -- CP-element group 1112: successors 
    -- CP-element group 1112: 	1115 
    -- CP-element group 1112:  members (1) 
      -- CP-element group 1112: 	 branch_block_stmt_714/merge_stmt_4132_PhiAck/phi_stmt_4133_ack
      -- 
    phi_stmt_4133_ack_13449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4133_ack_0, ack => zeropad3D_CP_2152_elements(1112)); -- 
    -- CP-element group 1113:  transition  input  bypass 
    -- CP-element group 1113: predecessors 
    -- CP-element group 1113: 	1111 
    -- CP-element group 1113: successors 
    -- CP-element group 1113: 	1115 
    -- CP-element group 1113:  members (1) 
      -- CP-element group 1113: 	 branch_block_stmt_714/merge_stmt_4132_PhiAck/phi_stmt_4140_ack
      -- 
    phi_stmt_4140_ack_13450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4140_ack_0, ack => zeropad3D_CP_2152_elements(1113)); -- 
    -- CP-element group 1114:  transition  input  bypass 
    -- CP-element group 1114: predecessors 
    -- CP-element group 1114: 	1111 
    -- CP-element group 1114: successors 
    -- CP-element group 1114: 	1115 
    -- CP-element group 1114:  members (1) 
      -- CP-element group 1114: 	 branch_block_stmt_714/merge_stmt_4132_PhiAck/phi_stmt_4146_ack
      -- 
    phi_stmt_4146_ack_13451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4146_ack_0, ack => zeropad3D_CP_2152_elements(1114)); -- 
    -- CP-element group 1115:  join  transition  bypass 
    -- CP-element group 1115: predecessors 
    -- CP-element group 1115: 	1112 
    -- CP-element group 1115: 	1113 
    -- CP-element group 1115: 	1114 
    -- CP-element group 1115: successors 
    -- CP-element group 1115: 	6 
    -- CP-element group 1115:  members (1) 
      -- CP-element group 1115: 	 branch_block_stmt_714/merge_stmt_4132_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1115: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1115"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1112) & zeropad3D_CP_2152_elements(1113) & zeropad3D_CP_2152_elements(1114);
      gj_zeropad3D_cp_element_group_1115 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1116:  transition  input  bypass 
    -- CP-element group 1116: predecessors 
    -- CP-element group 1116: 	592 
    -- CP-element group 1116: successors 
    -- CP-element group 1116: 	1118 
    -- CP-element group 1116:  members (2) 
      -- CP-element group 1116: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/type_cast_4158/SplitProtocol/Sample/$exit
      -- CP-element group 1116: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/type_cast_4158/SplitProtocol/Sample/ra
      -- 
    ra_13471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4158_inst_ack_0, ack => zeropad3D_CP_2152_elements(1116)); -- 
    -- CP-element group 1117:  transition  input  bypass 
    -- CP-element group 1117: predecessors 
    -- CP-element group 1117: 	592 
    -- CP-element group 1117: successors 
    -- CP-element group 1117: 	1118 
    -- CP-element group 1117:  members (2) 
      -- CP-element group 1117: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/type_cast_4158/SplitProtocol/Update/$exit
      -- CP-element group 1117: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/type_cast_4158/SplitProtocol/Update/ca
      -- 
    ca_13476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4158_inst_ack_1, ack => zeropad3D_CP_2152_elements(1117)); -- 
    -- CP-element group 1118:  join  transition  output  bypass 
    -- CP-element group 1118: predecessors 
    -- CP-element group 1118: 	1116 
    -- CP-element group 1118: 	1117 
    -- CP-element group 1118: successors 
    -- CP-element group 1118: 	1122 
    -- CP-element group 1118:  members (5) 
      -- CP-element group 1118: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/$exit
      -- CP-element group 1118: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/$exit
      -- CP-element group 1118: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/type_cast_4158/$exit
      -- CP-element group 1118: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_sources/type_cast_4158/SplitProtocol/$exit
      -- CP-element group 1118: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4155/phi_stmt_4155_req
      -- 
    phi_stmt_4155_req_13477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4155_req_13477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1118), ack => phi_stmt_4155_req_0); -- 
    zeropad3D_cp_element_group_1118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1116) & zeropad3D_CP_2152_elements(1117);
      gj_zeropad3D_cp_element_group_1118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1119:  transition  input  bypass 
    -- CP-element group 1119: predecessors 
    -- CP-element group 1119: 	592 
    -- CP-element group 1119: successors 
    -- CP-element group 1119: 	1121 
    -- CP-element group 1119:  members (2) 
      -- CP-element group 1119: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/type_cast_4162/SplitProtocol/Sample/$exit
      -- CP-element group 1119: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/type_cast_4162/SplitProtocol/Sample/ra
      -- 
    ra_13494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4162_inst_ack_0, ack => zeropad3D_CP_2152_elements(1119)); -- 
    -- CP-element group 1120:  transition  input  bypass 
    -- CP-element group 1120: predecessors 
    -- CP-element group 1120: 	592 
    -- CP-element group 1120: successors 
    -- CP-element group 1120: 	1121 
    -- CP-element group 1120:  members (2) 
      -- CP-element group 1120: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/type_cast_4162/SplitProtocol/Update/$exit
      -- CP-element group 1120: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/type_cast_4162/SplitProtocol/Update/ca
      -- 
    ca_13499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4162_inst_ack_1, ack => zeropad3D_CP_2152_elements(1120)); -- 
    -- CP-element group 1121:  join  transition  output  bypass 
    -- CP-element group 1121: predecessors 
    -- CP-element group 1121: 	1119 
    -- CP-element group 1121: 	1120 
    -- CP-element group 1121: successors 
    -- CP-element group 1121: 	1122 
    -- CP-element group 1121:  members (5) 
      -- CP-element group 1121: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/$exit
      -- CP-element group 1121: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/$exit
      -- CP-element group 1121: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/type_cast_4162/$exit
      -- CP-element group 1121: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_sources/type_cast_4162/SplitProtocol/$exit
      -- CP-element group 1121: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/phi_stmt_4159/phi_stmt_4159_req
      -- 
    phi_stmt_4159_req_13500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4159_req_13500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1121), ack => phi_stmt_4159_req_0); -- 
    zeropad3D_cp_element_group_1121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1119) & zeropad3D_CP_2152_elements(1120);
      gj_zeropad3D_cp_element_group_1121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1122:  join  fork  transition  place  bypass 
    -- CP-element group 1122: predecessors 
    -- CP-element group 1122: 	1118 
    -- CP-element group 1122: 	1121 
    -- CP-element group 1122: successors 
    -- CP-element group 1122: 	1123 
    -- CP-element group 1122: 	1124 
    -- CP-element group 1122:  members (3) 
      -- CP-element group 1122: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/$exit
      -- CP-element group 1122: 	 branch_block_stmt_714/merge_stmt_4154_PhiReqMerge
      -- CP-element group 1122: 	 branch_block_stmt_714/merge_stmt_4154_PhiAck/$entry
      -- 
    zeropad3D_cp_element_group_1122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1118) & zeropad3D_CP_2152_elements(1121);
      gj_zeropad3D_cp_element_group_1122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1123:  transition  input  bypass 
    -- CP-element group 1123: predecessors 
    -- CP-element group 1123: 	1122 
    -- CP-element group 1123: successors 
    -- CP-element group 1123: 	1125 
    -- CP-element group 1123:  members (1) 
      -- CP-element group 1123: 	 branch_block_stmt_714/merge_stmt_4154_PhiAck/phi_stmt_4155_ack
      -- 
    phi_stmt_4155_ack_13505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4155_ack_0, ack => zeropad3D_CP_2152_elements(1123)); -- 
    -- CP-element group 1124:  transition  input  bypass 
    -- CP-element group 1124: predecessors 
    -- CP-element group 1124: 	1122 
    -- CP-element group 1124: successors 
    -- CP-element group 1124: 	1125 
    -- CP-element group 1124:  members (1) 
      -- CP-element group 1124: 	 branch_block_stmt_714/merge_stmt_4154_PhiAck/phi_stmt_4159_ack
      -- 
    phi_stmt_4159_ack_13506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4159_ack_0, ack => zeropad3D_CP_2152_elements(1124)); -- 
    -- CP-element group 1125:  join  fork  transition  place  output  bypass 
    -- CP-element group 1125: predecessors 
    -- CP-element group 1125: 	1123 
    -- CP-element group 1125: 	1124 
    -- CP-element group 1125: successors 
    -- CP-element group 1125: 	594 
    -- CP-element group 1125: 	595 
    -- CP-element group 1125: 	596 
    -- CP-element group 1125: 	597 
    -- CP-element group 1125: 	598 
    -- CP-element group 1125: 	599 
    -- CP-element group 1125: 	600 
    -- CP-element group 1125: 	601 
    -- CP-element group 1125: 	602 
    -- CP-element group 1125: 	603 
    -- CP-element group 1125: 	605 
    -- CP-element group 1125: 	607 
    -- CP-element group 1125:  members (92) 
      -- CP-element group 1125: 	 branch_block_stmt_714/merge_stmt_4154__exit__
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293__entry__
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_update_start_
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_base_address_calculated
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_word_addrgen/root_register_ack
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_word_address_calculated
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Sample/word_access_start/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_root_address_calculated
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_base_address_resized
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_word_addrgen/root_register_req
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_sample_start_
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Update/word_access_complete/word_0/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Update/word_access_complete/word_0/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_word_addrgen/$exit
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Update/word_access_complete/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Update/word_access_complete/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_word_addrgen/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Update/word_access_complete/word_0/cr
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Update/word_access_complete/word_0/cr
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_base_plus_offset/sum_rename_ack
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Sample/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_base_plus_offset/sum_rename_req
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Update/word_access_complete/word_0/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Update/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Update/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Update/word_access_complete/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_base_plus_offset/$exit
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Sample/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Update/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Sample/word_access_start/word_0/rr
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Sample/word_access_start/word_0/rr
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Sample/word_access_start/word_0/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Sample/word_access_start/word_0/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Sample/word_access_start/word_0/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_root_address_calculated
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_word_address_calculated
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_update_start_
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_Sample/word_access_start/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Sample/word_access_start/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_sample_start_
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4166_Update/cr
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4166_Update/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_root_address_calculated
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_base_plus_offset/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_base_addr_resize/base_resize_ack
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_base_addr_resize/base_resize_req
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_base_addr_resize/$exit
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_word_address_calculated
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Sample/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4166_Sample/rr
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4166_Sample/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4166_update_start_
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4166_sample_start_
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_update_start_
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_base_addr_resize/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_depth_high_4184_sample_start_
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/LOAD_pad_4181_Sample/word_access_start/word_0/rr
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4196_Update/word_access_complete/word_0/cr
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_sample_start_
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_update_start_
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_base_address_calculated
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_word_address_calculated
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_root_address_calculated
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_base_address_resized
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_base_addr_resize/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_base_addr_resize/$exit
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_base_addr_resize/base_resize_req
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_base_addr_resize/base_resize_ack
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_base_plus_offset/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_base_plus_offset/$exit
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_base_plus_offset/sum_rename_req
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_base_plus_offset/sum_rename_ack
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_word_addrgen/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_word_addrgen/$exit
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_word_addrgen/root_register_req
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_word_addrgen/root_register_ack
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Sample/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Sample/word_access_start/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Sample/word_access_start/word_0/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Sample/word_access_start/word_0/rr
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Update/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Update/word_access_complete/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Update/word_access_complete/word_0/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/ptr_deref_4208_Update/word_access_complete/word_0/cr
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4212_update_start_
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4212_Update/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4212_Update/cr
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4251_update_start_
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4251_Update/$entry
      -- CP-element group 1125: 	 branch_block_stmt_714/assign_stmt_4167_to_assign_stmt_4293/type_cast_4251_Update/cr
      -- CP-element group 1125: 	 branch_block_stmt_714/merge_stmt_4154_PhiAck/$exit
      -- 
    cr_8992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1125), ack => LOAD_pad_4181_load_0_req_1); -- 
    cr_9025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1125), ack => LOAD_depth_high_4184_load_0_req_1); -- 
    rr_9014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1125), ack => LOAD_depth_high_4184_load_0_req_0); -- 
    rr_9064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1125), ack => ptr_deref_4196_load_0_req_0); -- 
    cr_8964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1125), ack => type_cast_4166_inst_req_1); -- 
    rr_8959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1125), ack => type_cast_4166_inst_req_0); -- 
    rr_8981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1125), ack => LOAD_pad_4181_load_0_req_0); -- 
    cr_9075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1125), ack => ptr_deref_4196_load_0_req_1); -- 
    rr_9114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1125), ack => ptr_deref_4208_load_0_req_0); -- 
    cr_9125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1125), ack => ptr_deref_4208_load_0_req_1); -- 
    cr_9144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1125), ack => type_cast_4212_inst_req_1); -- 
    cr_9158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1125), ack => type_cast_4251_inst_req_1); -- 
    zeropad3D_cp_element_group_1125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1123) & zeropad3D_CP_2152_elements(1124);
      gj_zeropad3D_cp_element_group_1125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1126:  transition  input  bypass 
    -- CP-element group 1126: predecessors 
    -- CP-element group 1126: 	7 
    -- CP-element group 1126: successors 
    -- CP-element group 1126: 	1128 
    -- CP-element group 1126:  members (2) 
      -- CP-element group 1126: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/type_cast_4302/SplitProtocol/Sample/$exit
      -- CP-element group 1126: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/type_cast_4302/SplitProtocol/Sample/ra
      -- 
    ra_13526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4302_inst_ack_0, ack => zeropad3D_CP_2152_elements(1126)); -- 
    -- CP-element group 1127:  transition  input  bypass 
    -- CP-element group 1127: predecessors 
    -- CP-element group 1127: 	7 
    -- CP-element group 1127: successors 
    -- CP-element group 1127: 	1128 
    -- CP-element group 1127:  members (2) 
      -- CP-element group 1127: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/type_cast_4302/SplitProtocol/Update/$exit
      -- CP-element group 1127: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/type_cast_4302/SplitProtocol/Update/ca
      -- 
    ca_13531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4302_inst_ack_1, ack => zeropad3D_CP_2152_elements(1127)); -- 
    -- CP-element group 1128:  join  transition  output  bypass 
    -- CP-element group 1128: predecessors 
    -- CP-element group 1128: 	1126 
    -- CP-element group 1128: 	1127 
    -- CP-element group 1128: successors 
    -- CP-element group 1128: 	1135 
    -- CP-element group 1128:  members (5) 
      -- CP-element group 1128: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/$exit
      -- CP-element group 1128: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/$exit
      -- CP-element group 1128: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/type_cast_4302/$exit
      -- CP-element group 1128: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/type_cast_4302/SplitProtocol/$exit
      -- CP-element group 1128: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_req
      -- 
    phi_stmt_4296_req_13532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4296_req_13532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1128), ack => phi_stmt_4296_req_1); -- 
    zeropad3D_cp_element_group_1128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1126) & zeropad3D_CP_2152_elements(1127);
      gj_zeropad3D_cp_element_group_1128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1129:  transition  input  bypass 
    -- CP-element group 1129: predecessors 
    -- CP-element group 1129: 	7 
    -- CP-element group 1129: successors 
    -- CP-element group 1129: 	1131 
    -- CP-element group 1129:  members (2) 
      -- CP-element group 1129: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4308/SplitProtocol/Sample/$exit
      -- CP-element group 1129: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4308/SplitProtocol/Sample/ra
      -- 
    ra_13549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4308_inst_ack_0, ack => zeropad3D_CP_2152_elements(1129)); -- 
    -- CP-element group 1130:  transition  input  bypass 
    -- CP-element group 1130: predecessors 
    -- CP-element group 1130: 	7 
    -- CP-element group 1130: successors 
    -- CP-element group 1130: 	1131 
    -- CP-element group 1130:  members (2) 
      -- CP-element group 1130: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4308/SplitProtocol/Update/$exit
      -- CP-element group 1130: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4308/SplitProtocol/Update/ca
      -- 
    ca_13554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4308_inst_ack_1, ack => zeropad3D_CP_2152_elements(1130)); -- 
    -- CP-element group 1131:  join  transition  output  bypass 
    -- CP-element group 1131: predecessors 
    -- CP-element group 1131: 	1129 
    -- CP-element group 1131: 	1130 
    -- CP-element group 1131: successors 
    -- CP-element group 1131: 	1135 
    -- CP-element group 1131:  members (5) 
      -- CP-element group 1131: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/$exit
      -- CP-element group 1131: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/$exit
      -- CP-element group 1131: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4308/$exit
      -- CP-element group 1131: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4308/SplitProtocol/$exit
      -- CP-element group 1131: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_req
      -- 
    phi_stmt_4303_req_13555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4303_req_13555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1131), ack => phi_stmt_4303_req_1); -- 
    zeropad3D_cp_element_group_1131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1129) & zeropad3D_CP_2152_elements(1130);
      gj_zeropad3D_cp_element_group_1131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1132:  transition  input  bypass 
    -- CP-element group 1132: predecessors 
    -- CP-element group 1132: 	7 
    -- CP-element group 1132: successors 
    -- CP-element group 1132: 	1134 
    -- CP-element group 1132:  members (2) 
      -- CP-element group 1132: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/type_cast_4315/SplitProtocol/Sample/$exit
      -- CP-element group 1132: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/type_cast_4315/SplitProtocol/Sample/ra
      -- 
    ra_13572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4315_inst_ack_0, ack => zeropad3D_CP_2152_elements(1132)); -- 
    -- CP-element group 1133:  transition  input  bypass 
    -- CP-element group 1133: predecessors 
    -- CP-element group 1133: 	7 
    -- CP-element group 1133: successors 
    -- CP-element group 1133: 	1134 
    -- CP-element group 1133:  members (2) 
      -- CP-element group 1133: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/type_cast_4315/SplitProtocol/Update/$exit
      -- CP-element group 1133: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/type_cast_4315/SplitProtocol/Update/ca
      -- 
    ca_13577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4315_inst_ack_1, ack => zeropad3D_CP_2152_elements(1133)); -- 
    -- CP-element group 1134:  join  transition  output  bypass 
    -- CP-element group 1134: predecessors 
    -- CP-element group 1134: 	1132 
    -- CP-element group 1134: 	1133 
    -- CP-element group 1134: successors 
    -- CP-element group 1134: 	1135 
    -- CP-element group 1134:  members (5) 
      -- CP-element group 1134: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/$exit
      -- CP-element group 1134: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/$exit
      -- CP-element group 1134: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/type_cast_4315/$exit
      -- CP-element group 1134: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/type_cast_4315/SplitProtocol/$exit
      -- CP-element group 1134: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_req
      -- 
    phi_stmt_4309_req_13578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4309_req_13578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1134), ack => phi_stmt_4309_req_1); -- 
    zeropad3D_cp_element_group_1134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1132) & zeropad3D_CP_2152_elements(1133);
      gj_zeropad3D_cp_element_group_1134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1135:  join  transition  bypass 
    -- CP-element group 1135: predecessors 
    -- CP-element group 1135: 	1128 
    -- CP-element group 1135: 	1131 
    -- CP-element group 1135: 	1134 
    -- CP-element group 1135: successors 
    -- CP-element group 1135: 	1142 
    -- CP-element group 1135:  members (1) 
      -- CP-element group 1135: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1135: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1135"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1128) & zeropad3D_CP_2152_elements(1131) & zeropad3D_CP_2152_elements(1134);
      gj_zeropad3D_cp_element_group_1135 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1136:  transition  output  delay-element  bypass 
    -- CP-element group 1136: predecessors 
    -- CP-element group 1136: 	608 
    -- CP-element group 1136: successors 
    -- CP-element group 1136: 	1141 
    -- CP-element group 1136:  members (4) 
      -- CP-element group 1136: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4296/$exit
      -- CP-element group 1136: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/$exit
      -- CP-element group 1136: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_sources/type_cast_4300_konst_delay_trans
      -- CP-element group 1136: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4296/phi_stmt_4296_req
      -- 
    phi_stmt_4296_req_13589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4296_req_13589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1136), ack => phi_stmt_4296_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(1136) is a control-delay.
    cp_element_1136_delay: control_delay_element  generic map(name => " 1136_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(608), ack => zeropad3D_CP_2152_elements(1136), clk => clk, reset =>reset);
    -- CP-element group 1137:  transition  input  bypass 
    -- CP-element group 1137: predecessors 
    -- CP-element group 1137: 	608 
    -- CP-element group 1137: successors 
    -- CP-element group 1137: 	1139 
    -- CP-element group 1137:  members (2) 
      -- CP-element group 1137: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4306/SplitProtocol/Sample/$exit
      -- CP-element group 1137: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4306/SplitProtocol/Sample/ra
      -- 
    ra_13606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4306_inst_ack_0, ack => zeropad3D_CP_2152_elements(1137)); -- 
    -- CP-element group 1138:  transition  input  bypass 
    -- CP-element group 1138: predecessors 
    -- CP-element group 1138: 	608 
    -- CP-element group 1138: successors 
    -- CP-element group 1138: 	1139 
    -- CP-element group 1138:  members (2) 
      -- CP-element group 1138: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4306/SplitProtocol/Update/$exit
      -- CP-element group 1138: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4306/SplitProtocol/Update/ca
      -- 
    ca_13611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4306_inst_ack_1, ack => zeropad3D_CP_2152_elements(1138)); -- 
    -- CP-element group 1139:  join  transition  output  bypass 
    -- CP-element group 1139: predecessors 
    -- CP-element group 1139: 	1137 
    -- CP-element group 1139: 	1138 
    -- CP-element group 1139: successors 
    -- CP-element group 1139: 	1141 
    -- CP-element group 1139:  members (5) 
      -- CP-element group 1139: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/$exit
      -- CP-element group 1139: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/$exit
      -- CP-element group 1139: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4306/$exit
      -- CP-element group 1139: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_sources/type_cast_4306/SplitProtocol/$exit
      -- CP-element group 1139: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4303/phi_stmt_4303_req
      -- 
    phi_stmt_4303_req_13612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4303_req_13612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1139), ack => phi_stmt_4303_req_0); -- 
    zeropad3D_cp_element_group_1139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1137) & zeropad3D_CP_2152_elements(1138);
      gj_zeropad3D_cp_element_group_1139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1140:  transition  output  delay-element  bypass 
    -- CP-element group 1140: predecessors 
    -- CP-element group 1140: 	608 
    -- CP-element group 1140: successors 
    -- CP-element group 1140: 	1141 
    -- CP-element group 1140:  members (4) 
      -- CP-element group 1140: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4309/$exit
      -- CP-element group 1140: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/$exit
      -- CP-element group 1140: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_sources/type_cast_4313_konst_delay_trans
      -- CP-element group 1140: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4309/phi_stmt_4309_req
      -- 
    phi_stmt_4309_req_13620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4309_req_13620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1140), ack => phi_stmt_4309_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(1140) is a control-delay.
    cp_element_1140_delay: control_delay_element  generic map(name => " 1140_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(608), ack => zeropad3D_CP_2152_elements(1140), clk => clk, reset =>reset);
    -- CP-element group 1141:  join  transition  bypass 
    -- CP-element group 1141: predecessors 
    -- CP-element group 1141: 	1136 
    -- CP-element group 1141: 	1139 
    -- CP-element group 1141: 	1140 
    -- CP-element group 1141: successors 
    -- CP-element group 1141: 	1142 
    -- CP-element group 1141:  members (1) 
      -- CP-element group 1141: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1141: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1141"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1136) & zeropad3D_CP_2152_elements(1139) & zeropad3D_CP_2152_elements(1140);
      gj_zeropad3D_cp_element_group_1141 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1142:  merge  fork  transition  place  bypass 
    -- CP-element group 1142: predecessors 
    -- CP-element group 1142: 	1135 
    -- CP-element group 1142: 	1141 
    -- CP-element group 1142: successors 
    -- CP-element group 1142: 	1143 
    -- CP-element group 1142: 	1144 
    -- CP-element group 1142: 	1145 
    -- CP-element group 1142:  members (2) 
      -- CP-element group 1142: 	 branch_block_stmt_714/merge_stmt_4295_PhiReqMerge
      -- CP-element group 1142: 	 branch_block_stmt_714/merge_stmt_4295_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1142) <= OrReduce(zeropad3D_CP_2152_elements(1135) & zeropad3D_CP_2152_elements(1141));
    -- CP-element group 1143:  transition  input  bypass 
    -- CP-element group 1143: predecessors 
    -- CP-element group 1143: 	1142 
    -- CP-element group 1143: successors 
    -- CP-element group 1143: 	1146 
    -- CP-element group 1143:  members (1) 
      -- CP-element group 1143: 	 branch_block_stmt_714/merge_stmt_4295_PhiAck/phi_stmt_4296_ack
      -- 
    phi_stmt_4296_ack_13625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4296_ack_0, ack => zeropad3D_CP_2152_elements(1143)); -- 
    -- CP-element group 1144:  transition  input  bypass 
    -- CP-element group 1144: predecessors 
    -- CP-element group 1144: 	1142 
    -- CP-element group 1144: successors 
    -- CP-element group 1144: 	1146 
    -- CP-element group 1144:  members (1) 
      -- CP-element group 1144: 	 branch_block_stmt_714/merge_stmt_4295_PhiAck/phi_stmt_4303_ack
      -- 
    phi_stmt_4303_ack_13626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4303_ack_0, ack => zeropad3D_CP_2152_elements(1144)); -- 
    -- CP-element group 1145:  transition  input  bypass 
    -- CP-element group 1145: predecessors 
    -- CP-element group 1145: 	1142 
    -- CP-element group 1145: successors 
    -- CP-element group 1145: 	1146 
    -- CP-element group 1145:  members (1) 
      -- CP-element group 1145: 	 branch_block_stmt_714/merge_stmt_4295_PhiAck/phi_stmt_4309_ack
      -- 
    phi_stmt_4309_ack_13627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4309_ack_0, ack => zeropad3D_CP_2152_elements(1145)); -- 
    -- CP-element group 1146:  join  fork  transition  place  output  bypass 
    -- CP-element group 1146: predecessors 
    -- CP-element group 1146: 	1143 
    -- CP-element group 1146: 	1144 
    -- CP-element group 1146: 	1145 
    -- CP-element group 1146: successors 
    -- CP-element group 1146: 	609 
    -- CP-element group 1146: 	610 
    -- CP-element group 1146:  members (10) 
      -- CP-element group 1146: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328__entry__
      -- CP-element group 1146: 	 branch_block_stmt_714/merge_stmt_4295__exit__
      -- CP-element group 1146: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/$entry
      -- CP-element group 1146: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/type_cast_4320_sample_start_
      -- CP-element group 1146: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/type_cast_4320_update_start_
      -- CP-element group 1146: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/type_cast_4320_Sample/$entry
      -- CP-element group 1146: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/type_cast_4320_Sample/rr
      -- CP-element group 1146: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/type_cast_4320_Update/$entry
      -- CP-element group 1146: 	 branch_block_stmt_714/assign_stmt_4321_to_assign_stmt_4328/type_cast_4320_Update/cr
      -- CP-element group 1146: 	 branch_block_stmt_714/merge_stmt_4295_PhiAck/$exit
      -- 
    rr_9170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1146), ack => type_cast_4320_inst_req_0); -- 
    cr_9175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1146), ack => type_cast_4320_inst_req_1); -- 
    zeropad3D_cp_element_group_1146: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1146"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1143) & zeropad3D_CP_2152_elements(1144) & zeropad3D_CP_2152_elements(1145);
      gj_zeropad3D_cp_element_group_1146 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1147:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1147: predecessors 
    -- CP-element group 1147: 	611 
    -- CP-element group 1147: 	618 
    -- CP-element group 1147: 	621 
    -- CP-element group 1147: 	628 
    -- CP-element group 1147: successors 
    -- CP-element group 1147: 	629 
    -- CP-element group 1147: 	630 
    -- CP-element group 1147: 	631 
    -- CP-element group 1147: 	632 
    -- CP-element group 1147: 	635 
    -- CP-element group 1147: 	637 
    -- CP-element group 1147: 	639 
    -- CP-element group 1147: 	641 
    -- CP-element group 1147:  members (33) 
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468__entry__
      -- CP-element group 1147: 	 branch_block_stmt_714/merge_stmt_4412__exit__
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/$entry
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4416_sample_start_
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4416_update_start_
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4416_Sample/$entry
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4416_Sample/rr
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4416_Update/$entry
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4416_Update/cr
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4421_sample_start_
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4421_update_start_
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4421_Sample/$entry
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4421_Sample/rr
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4421_Update/$entry
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4421_Update/cr
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4455_update_start_
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4455_Update/$entry
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/type_cast_4455_Update/cr
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/addr_of_4462_update_start_
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_final_index_sum_regn_update_start
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_final_index_sum_regn_Update/$entry
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/array_obj_ref_4461_final_index_sum_regn_Update/req
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/addr_of_4462_complete/$entry
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/addr_of_4462_complete/req
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_update_start_
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Update/$entry
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Update/word_access_complete/$entry
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Update/word_access_complete/word_0/$entry
      -- CP-element group 1147: 	 branch_block_stmt_714/assign_stmt_4417_to_assign_stmt_4468/ptr_deref_4465_Update/word_access_complete/word_0/cr
      -- CP-element group 1147: 	 branch_block_stmt_714/merge_stmt_4412_PhiReqMerge
      -- CP-element group 1147: 	 branch_block_stmt_714/merge_stmt_4412_PhiAck/$entry
      -- CP-element group 1147: 	 branch_block_stmt_714/merge_stmt_4412_PhiAck/$exit
      -- CP-element group 1147: 	 branch_block_stmt_714/merge_stmt_4412_PhiAck/dummy
      -- 
    rr_9380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1147), ack => type_cast_4416_inst_req_0); -- 
    cr_9385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1147), ack => type_cast_4416_inst_req_1); -- 
    rr_9394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1147), ack => type_cast_4421_inst_req_0); -- 
    cr_9399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1147), ack => type_cast_4421_inst_req_1); -- 
    cr_9413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1147), ack => type_cast_4455_inst_req_1); -- 
    req_9444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1147), ack => array_obj_ref_4461_index_offset_req_1); -- 
    req_9459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1147), ack => addr_of_4462_final_reg_req_1); -- 
    cr_9509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1147), ack => ptr_deref_4465_store_0_req_1); -- 
    zeropad3D_CP_2152_elements(1147) <= OrReduce(zeropad3D_CP_2152_elements(611) & zeropad3D_CP_2152_elements(618) & zeropad3D_CP_2152_elements(621) & zeropad3D_CP_2152_elements(628));
    -- CP-element group 1148:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1148: predecessors 
    -- CP-element group 1148: 	642 
    -- CP-element group 1148: 	662 
    -- CP-element group 1148: successors 
    -- CP-element group 1148: 	663 
    -- CP-element group 1148: 	664 
    -- CP-element group 1148:  members (13) 
      -- CP-element group 1148: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595__entry__
      -- CP-element group 1148: 	 branch_block_stmt_714/merge_stmt_4577__exit__
      -- CP-element group 1148: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/type_cast_4581_update_start_
      -- CP-element group 1148: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/type_cast_4581_sample_start_
      -- CP-element group 1148: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/type_cast_4581_Update/cr
      -- CP-element group 1148: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/$entry
      -- CP-element group 1148: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/type_cast_4581_Update/$entry
      -- CP-element group 1148: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/type_cast_4581_Sample/rr
      -- CP-element group 1148: 	 branch_block_stmt_714/assign_stmt_4582_to_assign_stmt_4595/type_cast_4581_Sample/$entry
      -- CP-element group 1148: 	 branch_block_stmt_714/merge_stmt_4577_PhiReqMerge
      -- CP-element group 1148: 	 branch_block_stmt_714/merge_stmt_4577_PhiAck/$entry
      -- CP-element group 1148: 	 branch_block_stmt_714/merge_stmt_4577_PhiAck/$exit
      -- CP-element group 1148: 	 branch_block_stmt_714/merge_stmt_4577_PhiAck/dummy
      -- 
    cr_9763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1148), ack => type_cast_4581_inst_req_1); -- 
    rr_9758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1148), ack => type_cast_4581_inst_req_0); -- 
    zeropad3D_CP_2152_elements(1148) <= OrReduce(zeropad3D_CP_2152_elements(642) & zeropad3D_CP_2152_elements(662));
    -- CP-element group 1149:  transition  input  bypass 
    -- CP-element group 1149: predecessors 
    -- CP-element group 1149: 	684 
    -- CP-element group 1149: successors 
    -- CP-element group 1149: 	1151 
    -- CP-element group 1149:  members (2) 
      -- CP-element group 1149: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4706/SplitProtocol/Sample/$exit
      -- CP-element group 1149: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4706/SplitProtocol/Sample/ra
      -- 
    ra_13747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4706_inst_ack_0, ack => zeropad3D_CP_2152_elements(1149)); -- 
    -- CP-element group 1150:  transition  input  bypass 
    -- CP-element group 1150: predecessors 
    -- CP-element group 1150: 	684 
    -- CP-element group 1150: successors 
    -- CP-element group 1150: 	1151 
    -- CP-element group 1150:  members (2) 
      -- CP-element group 1150: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4706/SplitProtocol/Update/$exit
      -- CP-element group 1150: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4706/SplitProtocol/Update/ca
      -- 
    ca_13752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4706_inst_ack_1, ack => zeropad3D_CP_2152_elements(1150)); -- 
    -- CP-element group 1151:  join  transition  output  bypass 
    -- CP-element group 1151: predecessors 
    -- CP-element group 1151: 	1149 
    -- CP-element group 1151: 	1150 
    -- CP-element group 1151: successors 
    -- CP-element group 1151: 	1156 
    -- CP-element group 1151:  members (5) 
      -- CP-element group 1151: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/$exit
      -- CP-element group 1151: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/$exit
      -- CP-element group 1151: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4706/$exit
      -- CP-element group 1151: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4706/SplitProtocol/$exit
      -- CP-element group 1151: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_req
      -- 
    phi_stmt_4703_req_13753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4703_req_13753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1151), ack => phi_stmt_4703_req_0); -- 
    zeropad3D_cp_element_group_1151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1149) & zeropad3D_CP_2152_elements(1150);
      gj_zeropad3D_cp_element_group_1151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1152:  transition  input  bypass 
    -- CP-element group 1152: predecessors 
    -- CP-element group 1152: 	684 
    -- CP-element group 1152: successors 
    -- CP-element group 1152: 	1154 
    -- CP-element group 1152:  members (2) 
      -- CP-element group 1152: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4702/SplitProtocol/Sample/$exit
      -- CP-element group 1152: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4702/SplitProtocol/Sample/ra
      -- 
    ra_13770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4702_inst_ack_0, ack => zeropad3D_CP_2152_elements(1152)); -- 
    -- CP-element group 1153:  transition  input  bypass 
    -- CP-element group 1153: predecessors 
    -- CP-element group 1153: 	684 
    -- CP-element group 1153: successors 
    -- CP-element group 1153: 	1154 
    -- CP-element group 1153:  members (2) 
      -- CP-element group 1153: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4702/SplitProtocol/Update/$exit
      -- CP-element group 1153: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4702/SplitProtocol/Update/ca
      -- 
    ca_13775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4702_inst_ack_1, ack => zeropad3D_CP_2152_elements(1153)); -- 
    -- CP-element group 1154:  join  transition  output  bypass 
    -- CP-element group 1154: predecessors 
    -- CP-element group 1154: 	1152 
    -- CP-element group 1154: 	1153 
    -- CP-element group 1154: successors 
    -- CP-element group 1154: 	1156 
    -- CP-element group 1154:  members (5) 
      -- CP-element group 1154: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/$exit
      -- CP-element group 1154: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/$exit
      -- CP-element group 1154: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4702/$exit
      -- CP-element group 1154: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4702/SplitProtocol/$exit
      -- CP-element group 1154: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_req
      -- 
    phi_stmt_4697_req_13776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4697_req_13776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1154), ack => phi_stmt_4697_req_1); -- 
    zeropad3D_cp_element_group_1154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1152) & zeropad3D_CP_2152_elements(1153);
      gj_zeropad3D_cp_element_group_1154 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1155:  transition  output  delay-element  bypass 
    -- CP-element group 1155: predecessors 
    -- CP-element group 1155: 	684 
    -- CP-element group 1155: successors 
    -- CP-element group 1155: 	1156 
    -- CP-element group 1155:  members (4) 
      -- CP-element group 1155: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4690/$exit
      -- CP-element group 1155: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/$exit
      -- CP-element group 1155: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/type_cast_4694_konst_delay_trans
      -- CP-element group 1155: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_req
      -- 
    phi_stmt_4690_req_13784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4690_req_13784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1155), ack => phi_stmt_4690_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(1155) is a control-delay.
    cp_element_1155_delay: control_delay_element  generic map(name => " 1155_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(684), ack => zeropad3D_CP_2152_elements(1155), clk => clk, reset =>reset);
    -- CP-element group 1156:  join  transition  bypass 
    -- CP-element group 1156: predecessors 
    -- CP-element group 1156: 	1151 
    -- CP-element group 1156: 	1154 
    -- CP-element group 1156: 	1155 
    -- CP-element group 1156: successors 
    -- CP-element group 1156: 	1167 
    -- CP-element group 1156:  members (1) 
      -- CP-element group 1156: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1156: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1156"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1151) & zeropad3D_CP_2152_elements(1154) & zeropad3D_CP_2152_elements(1155);
      gj_zeropad3D_cp_element_group_1156 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1157:  transition  input  bypass 
    -- CP-element group 1157: predecessors 
    -- CP-element group 1157: 	665 
    -- CP-element group 1157: successors 
    -- CP-element group 1157: 	1159 
    -- CP-element group 1157:  members (2) 
      -- CP-element group 1157: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4708/SplitProtocol/Sample/$exit
      -- CP-element group 1157: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4708/SplitProtocol/Sample/ra
      -- 
    ra_13804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4708_inst_ack_0, ack => zeropad3D_CP_2152_elements(1157)); -- 
    -- CP-element group 1158:  transition  input  bypass 
    -- CP-element group 1158: predecessors 
    -- CP-element group 1158: 	665 
    -- CP-element group 1158: successors 
    -- CP-element group 1158: 	1159 
    -- CP-element group 1158:  members (2) 
      -- CP-element group 1158: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4708/SplitProtocol/Update/$exit
      -- CP-element group 1158: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4708/SplitProtocol/Update/ca
      -- 
    ca_13809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4708_inst_ack_1, ack => zeropad3D_CP_2152_elements(1158)); -- 
    -- CP-element group 1159:  join  transition  output  bypass 
    -- CP-element group 1159: predecessors 
    -- CP-element group 1159: 	1157 
    -- CP-element group 1159: 	1158 
    -- CP-element group 1159: successors 
    -- CP-element group 1159: 	1166 
    -- CP-element group 1159:  members (5) 
      -- CP-element group 1159: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/$exit
      -- CP-element group 1159: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/$exit
      -- CP-element group 1159: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4708/$exit
      -- CP-element group 1159: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_sources/type_cast_4708/SplitProtocol/$exit
      -- CP-element group 1159: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4703/phi_stmt_4703_req
      -- 
    phi_stmt_4703_req_13810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4703_req_13810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1159), ack => phi_stmt_4703_req_1); -- 
    zeropad3D_cp_element_group_1159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1157) & zeropad3D_CP_2152_elements(1158);
      gj_zeropad3D_cp_element_group_1159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1160:  transition  input  bypass 
    -- CP-element group 1160: predecessors 
    -- CP-element group 1160: 	665 
    -- CP-element group 1160: successors 
    -- CP-element group 1160: 	1162 
    -- CP-element group 1160:  members (2) 
      -- CP-element group 1160: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4700/SplitProtocol/Sample/$exit
      -- CP-element group 1160: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4700/SplitProtocol/Sample/ra
      -- 
    ra_13827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4700_inst_ack_0, ack => zeropad3D_CP_2152_elements(1160)); -- 
    -- CP-element group 1161:  transition  input  bypass 
    -- CP-element group 1161: predecessors 
    -- CP-element group 1161: 	665 
    -- CP-element group 1161: successors 
    -- CP-element group 1161: 	1162 
    -- CP-element group 1161:  members (2) 
      -- CP-element group 1161: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4700/SplitProtocol/Update/$exit
      -- CP-element group 1161: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4700/SplitProtocol/Update/ca
      -- 
    ca_13832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4700_inst_ack_1, ack => zeropad3D_CP_2152_elements(1161)); -- 
    -- CP-element group 1162:  join  transition  output  bypass 
    -- CP-element group 1162: predecessors 
    -- CP-element group 1162: 	1160 
    -- CP-element group 1162: 	1161 
    -- CP-element group 1162: successors 
    -- CP-element group 1162: 	1166 
    -- CP-element group 1162:  members (5) 
      -- CP-element group 1162: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/$exit
      -- CP-element group 1162: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/$exit
      -- CP-element group 1162: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4700/$exit
      -- CP-element group 1162: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_sources/type_cast_4700/SplitProtocol/$exit
      -- CP-element group 1162: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4697/phi_stmt_4697_req
      -- 
    phi_stmt_4697_req_13833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4697_req_13833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1162), ack => phi_stmt_4697_req_0); -- 
    zeropad3D_cp_element_group_1162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1160) & zeropad3D_CP_2152_elements(1161);
      gj_zeropad3D_cp_element_group_1162 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1163:  transition  input  bypass 
    -- CP-element group 1163: predecessors 
    -- CP-element group 1163: 	665 
    -- CP-element group 1163: successors 
    -- CP-element group 1163: 	1165 
    -- CP-element group 1163:  members (2) 
      -- CP-element group 1163: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/type_cast_4696/SplitProtocol/Sample/$exit
      -- CP-element group 1163: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/type_cast_4696/SplitProtocol/Sample/ra
      -- 
    ra_13850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4696_inst_ack_0, ack => zeropad3D_CP_2152_elements(1163)); -- 
    -- CP-element group 1164:  transition  input  bypass 
    -- CP-element group 1164: predecessors 
    -- CP-element group 1164: 	665 
    -- CP-element group 1164: successors 
    -- CP-element group 1164: 	1165 
    -- CP-element group 1164:  members (2) 
      -- CP-element group 1164: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/type_cast_4696/SplitProtocol/Update/$exit
      -- CP-element group 1164: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/type_cast_4696/SplitProtocol/Update/ca
      -- 
    ca_13855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4696_inst_ack_1, ack => zeropad3D_CP_2152_elements(1164)); -- 
    -- CP-element group 1165:  join  transition  output  bypass 
    -- CP-element group 1165: predecessors 
    -- CP-element group 1165: 	1163 
    -- CP-element group 1165: 	1164 
    -- CP-element group 1165: successors 
    -- CP-element group 1165: 	1166 
    -- CP-element group 1165:  members (5) 
      -- CP-element group 1165: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/$exit
      -- CP-element group 1165: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/$exit
      -- CP-element group 1165: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/type_cast_4696/$exit
      -- CP-element group 1165: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_sources/type_cast_4696/SplitProtocol/$exit
      -- CP-element group 1165: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4690/phi_stmt_4690_req
      -- 
    phi_stmt_4690_req_13856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4690_req_13856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1165), ack => phi_stmt_4690_req_1); -- 
    zeropad3D_cp_element_group_1165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1163) & zeropad3D_CP_2152_elements(1164);
      gj_zeropad3D_cp_element_group_1165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1166:  join  transition  bypass 
    -- CP-element group 1166: predecessors 
    -- CP-element group 1166: 	1159 
    -- CP-element group 1166: 	1162 
    -- CP-element group 1166: 	1165 
    -- CP-element group 1166: successors 
    -- CP-element group 1166: 	1167 
    -- CP-element group 1166:  members (1) 
      -- CP-element group 1166: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1166: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1166"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1159) & zeropad3D_CP_2152_elements(1162) & zeropad3D_CP_2152_elements(1165);
      gj_zeropad3D_cp_element_group_1166 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1167:  merge  fork  transition  place  bypass 
    -- CP-element group 1167: predecessors 
    -- CP-element group 1167: 	1156 
    -- CP-element group 1167: 	1166 
    -- CP-element group 1167: successors 
    -- CP-element group 1167: 	1168 
    -- CP-element group 1167: 	1169 
    -- CP-element group 1167: 	1170 
    -- CP-element group 1167:  members (2) 
      -- CP-element group 1167: 	 branch_block_stmt_714/merge_stmt_4689_PhiReqMerge
      -- CP-element group 1167: 	 branch_block_stmt_714/merge_stmt_4689_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1167) <= OrReduce(zeropad3D_CP_2152_elements(1156) & zeropad3D_CP_2152_elements(1166));
    -- CP-element group 1168:  transition  input  bypass 
    -- CP-element group 1168: predecessors 
    -- CP-element group 1168: 	1167 
    -- CP-element group 1168: successors 
    -- CP-element group 1168: 	1171 
    -- CP-element group 1168:  members (1) 
      -- CP-element group 1168: 	 branch_block_stmt_714/merge_stmt_4689_PhiAck/phi_stmt_4690_ack
      -- 
    phi_stmt_4690_ack_13861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4690_ack_0, ack => zeropad3D_CP_2152_elements(1168)); -- 
    -- CP-element group 1169:  transition  input  bypass 
    -- CP-element group 1169: predecessors 
    -- CP-element group 1169: 	1167 
    -- CP-element group 1169: successors 
    -- CP-element group 1169: 	1171 
    -- CP-element group 1169:  members (1) 
      -- CP-element group 1169: 	 branch_block_stmt_714/merge_stmt_4689_PhiAck/phi_stmt_4697_ack
      -- 
    phi_stmt_4697_ack_13862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4697_ack_0, ack => zeropad3D_CP_2152_elements(1169)); -- 
    -- CP-element group 1170:  transition  input  bypass 
    -- CP-element group 1170: predecessors 
    -- CP-element group 1170: 	1167 
    -- CP-element group 1170: successors 
    -- CP-element group 1170: 	1171 
    -- CP-element group 1170:  members (1) 
      -- CP-element group 1170: 	 branch_block_stmt_714/merge_stmt_4689_PhiAck/phi_stmt_4703_ack
      -- 
    phi_stmt_4703_ack_13863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4703_ack_0, ack => zeropad3D_CP_2152_elements(1170)); -- 
    -- CP-element group 1171:  join  transition  bypass 
    -- CP-element group 1171: predecessors 
    -- CP-element group 1171: 	1168 
    -- CP-element group 1171: 	1169 
    -- CP-element group 1171: 	1170 
    -- CP-element group 1171: successors 
    -- CP-element group 1171: 	7 
    -- CP-element group 1171:  members (1) 
      -- CP-element group 1171: 	 branch_block_stmt_714/merge_stmt_4689_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1171: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1171"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1168) & zeropad3D_CP_2152_elements(1169) & zeropad3D_CP_2152_elements(1170);
      gj_zeropad3D_cp_element_group_1171 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1172:  transition  input  bypass 
    -- CP-element group 1172: predecessors 
    -- CP-element group 1172: 	683 
    -- CP-element group 1172: successors 
    -- CP-element group 1172: 	1174 
    -- CP-element group 1172:  members (2) 
      -- CP-element group 1172: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/type_cast_4719/SplitProtocol/Sample/$exit
      -- CP-element group 1172: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/type_cast_4719/SplitProtocol/Sample/ra
      -- 
    ra_13883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4719_inst_ack_0, ack => zeropad3D_CP_2152_elements(1172)); -- 
    -- CP-element group 1173:  transition  input  bypass 
    -- CP-element group 1173: predecessors 
    -- CP-element group 1173: 	683 
    -- CP-element group 1173: successors 
    -- CP-element group 1173: 	1174 
    -- CP-element group 1173:  members (2) 
      -- CP-element group 1173: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/type_cast_4719/SplitProtocol/Update/$exit
      -- CP-element group 1173: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/type_cast_4719/SplitProtocol/Update/ca
      -- 
    ca_13888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4719_inst_ack_1, ack => zeropad3D_CP_2152_elements(1173)); -- 
    -- CP-element group 1174:  join  transition  output  bypass 
    -- CP-element group 1174: predecessors 
    -- CP-element group 1174: 	1172 
    -- CP-element group 1174: 	1173 
    -- CP-element group 1174: successors 
    -- CP-element group 1174: 	1181 
    -- CP-element group 1174:  members (5) 
      -- CP-element group 1174: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/$exit
      -- CP-element group 1174: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/$exit
      -- CP-element group 1174: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/type_cast_4719/$exit
      -- CP-element group 1174: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_sources/type_cast_4719/SplitProtocol/$exit
      -- CP-element group 1174: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4716/phi_stmt_4716_req
      -- 
    phi_stmt_4716_req_13889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4716_req_13889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1174), ack => phi_stmt_4716_req_0); -- 
    zeropad3D_cp_element_group_1174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1172) & zeropad3D_CP_2152_elements(1173);
      gj_zeropad3D_cp_element_group_1174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1175:  transition  input  bypass 
    -- CP-element group 1175: predecessors 
    -- CP-element group 1175: 	683 
    -- CP-element group 1175: successors 
    -- CP-element group 1175: 	1177 
    -- CP-element group 1175:  members (2) 
      -- CP-element group 1175: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/type_cast_4715/SplitProtocol/Sample/$exit
      -- CP-element group 1175: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/type_cast_4715/SplitProtocol/Sample/ra
      -- 
    ra_13906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4715_inst_ack_0, ack => zeropad3D_CP_2152_elements(1175)); -- 
    -- CP-element group 1176:  transition  input  bypass 
    -- CP-element group 1176: predecessors 
    -- CP-element group 1176: 	683 
    -- CP-element group 1176: successors 
    -- CP-element group 1176: 	1177 
    -- CP-element group 1176:  members (2) 
      -- CP-element group 1176: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/type_cast_4715/SplitProtocol/Update/$exit
      -- CP-element group 1176: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/type_cast_4715/SplitProtocol/Update/ca
      -- 
    ca_13911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4715_inst_ack_1, ack => zeropad3D_CP_2152_elements(1176)); -- 
    -- CP-element group 1177:  join  transition  output  bypass 
    -- CP-element group 1177: predecessors 
    -- CP-element group 1177: 	1175 
    -- CP-element group 1177: 	1176 
    -- CP-element group 1177: successors 
    -- CP-element group 1177: 	1181 
    -- CP-element group 1177:  members (5) 
      -- CP-element group 1177: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/$exit
      -- CP-element group 1177: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/$exit
      -- CP-element group 1177: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/type_cast_4715/$exit
      -- CP-element group 1177: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_sources/type_cast_4715/SplitProtocol/$exit
      -- CP-element group 1177: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4712/phi_stmt_4712_req
      -- 
    phi_stmt_4712_req_13912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4712_req_13912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1177), ack => phi_stmt_4712_req_0); -- 
    zeropad3D_cp_element_group_1177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1175) & zeropad3D_CP_2152_elements(1176);
      gj_zeropad3D_cp_element_group_1177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1178:  transition  input  bypass 
    -- CP-element group 1178: predecessors 
    -- CP-element group 1178: 	683 
    -- CP-element group 1178: successors 
    -- CP-element group 1178: 	1180 
    -- CP-element group 1178:  members (2) 
      -- CP-element group 1178: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/type_cast_4723/SplitProtocol/Sample/$exit
      -- CP-element group 1178: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/type_cast_4723/SplitProtocol/Sample/ra
      -- 
    ra_13929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4723_inst_ack_0, ack => zeropad3D_CP_2152_elements(1178)); -- 
    -- CP-element group 1179:  transition  input  bypass 
    -- CP-element group 1179: predecessors 
    -- CP-element group 1179: 	683 
    -- CP-element group 1179: successors 
    -- CP-element group 1179: 	1180 
    -- CP-element group 1179:  members (2) 
      -- CP-element group 1179: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/type_cast_4723/SplitProtocol/Update/$exit
      -- CP-element group 1179: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/type_cast_4723/SplitProtocol/Update/ca
      -- 
    ca_13934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4723_inst_ack_1, ack => zeropad3D_CP_2152_elements(1179)); -- 
    -- CP-element group 1180:  join  transition  output  bypass 
    -- CP-element group 1180: predecessors 
    -- CP-element group 1180: 	1178 
    -- CP-element group 1180: 	1179 
    -- CP-element group 1180: successors 
    -- CP-element group 1180: 	1181 
    -- CP-element group 1180:  members (5) 
      -- CP-element group 1180: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/$exit
      -- CP-element group 1180: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/$exit
      -- CP-element group 1180: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/type_cast_4723/$exit
      -- CP-element group 1180: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_sources/type_cast_4723/SplitProtocol/$exit
      -- CP-element group 1180: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/phi_stmt_4720/phi_stmt_4720_req
      -- 
    phi_stmt_4720_req_13935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4720_req_13935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1180), ack => phi_stmt_4720_req_0); -- 
    zeropad3D_cp_element_group_1180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1178) & zeropad3D_CP_2152_elements(1179);
      gj_zeropad3D_cp_element_group_1180 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1181:  join  fork  transition  place  bypass 
    -- CP-element group 1181: predecessors 
    -- CP-element group 1181: 	1174 
    -- CP-element group 1181: 	1177 
    -- CP-element group 1181: 	1180 
    -- CP-element group 1181: successors 
    -- CP-element group 1181: 	1182 
    -- CP-element group 1181: 	1183 
    -- CP-element group 1181: 	1184 
    -- CP-element group 1181:  members (3) 
      -- CP-element group 1181: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/$exit
      -- CP-element group 1181: 	 branch_block_stmt_714/merge_stmt_4711_PhiReqMerge
      -- CP-element group 1181: 	 branch_block_stmt_714/merge_stmt_4711_PhiAck/$entry
      -- 
    zeropad3D_cp_element_group_1181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1174) & zeropad3D_CP_2152_elements(1177) & zeropad3D_CP_2152_elements(1180);
      gj_zeropad3D_cp_element_group_1181 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1182:  transition  input  bypass 
    -- CP-element group 1182: predecessors 
    -- CP-element group 1182: 	1181 
    -- CP-element group 1182: successors 
    -- CP-element group 1182: 	1185 
    -- CP-element group 1182:  members (1) 
      -- CP-element group 1182: 	 branch_block_stmt_714/merge_stmt_4711_PhiAck/phi_stmt_4712_ack
      -- 
    phi_stmt_4712_ack_13940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4712_ack_0, ack => zeropad3D_CP_2152_elements(1182)); -- 
    -- CP-element group 1183:  transition  input  bypass 
    -- CP-element group 1183: predecessors 
    -- CP-element group 1183: 	1181 
    -- CP-element group 1183: successors 
    -- CP-element group 1183: 	1185 
    -- CP-element group 1183:  members (1) 
      -- CP-element group 1183: 	 branch_block_stmt_714/merge_stmt_4711_PhiAck/phi_stmt_4716_ack
      -- 
    phi_stmt_4716_ack_13941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4716_ack_0, ack => zeropad3D_CP_2152_elements(1183)); -- 
    -- CP-element group 1184:  transition  input  bypass 
    -- CP-element group 1184: predecessors 
    -- CP-element group 1184: 	1181 
    -- CP-element group 1184: successors 
    -- CP-element group 1184: 	1185 
    -- CP-element group 1184:  members (1) 
      -- CP-element group 1184: 	 branch_block_stmt_714/merge_stmt_4711_PhiAck/phi_stmt_4720_ack
      -- 
    phi_stmt_4720_ack_13942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4720_ack_0, ack => zeropad3D_CP_2152_elements(1184)); -- 
    -- CP-element group 1185:  join  fork  transition  place  output  bypass 
    -- CP-element group 1185: predecessors 
    -- CP-element group 1185: 	1182 
    -- CP-element group 1185: 	1183 
    -- CP-element group 1185: 	1184 
    -- CP-element group 1185: successors 
    -- CP-element group 1185: 	685 
    -- CP-element group 1185: 	686 
    -- CP-element group 1185: 	687 
    -- CP-element group 1185: 	688 
    -- CP-element group 1185: 	689 
    -- CP-element group 1185: 	690 
    -- CP-element group 1185: 	691 
    -- CP-element group 1185: 	692 
    -- CP-element group 1185: 	693 
    -- CP-element group 1185: 	694 
    -- CP-element group 1185: 	695 
    -- CP-element group 1185: 	696 
    -- CP-element group 1185: 	698 
    -- CP-element group 1185: 	700 
    -- CP-element group 1185:  members (98) 
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864__entry__
      -- CP-element group 1185: 	 branch_block_stmt_714/merge_stmt_4711__exit__
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Sample/word_access_start/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_base_plus_offset/sum_rename_req
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_base_plus_offset/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Sample/word_access_start/word_0/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_base_plus_offset/sum_rename_ack
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_base_plus_offset/$exit
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Sample/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_base_plus_offset/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_root_address_calculated
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_base_addr_resize/base_resize_ack
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_word_address_calculated
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_update_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_sample_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4737_Update/cr
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4783_Update/cr
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4737_Update/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_base_addr_resize/base_resize_ack
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Sample/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_base_addr_resize/base_resize_req
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Update/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_base_addr_resize/$exit
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_base_addr_resize/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4737_Sample/rr
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_base_address_resized
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4783_Update/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_root_address_calculated
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_word_address_calculated
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Sample/word_access_start/word_0/rr
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_word_addrgen/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_word_addrgen/root_register_ack
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_base_addr_resize/base_resize_req
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_base_address_calculated
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4737_Sample/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4737_update_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_base_addr_resize/$exit
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_base_addr_resize/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_base_address_resized
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_update_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_root_address_calculated
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4737_sample_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_sample_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4727_Update/cr
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_word_address_calculated
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_base_address_calculated
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_update_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_sample_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4727_Update/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Sample/word_access_start/word_0/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Sample/word_access_start/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4727_Sample/rr
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4727_Sample/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4822_Update/cr
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Update/word_access_complete/word_0/cr
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Update/word_access_complete/word_0/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4727_update_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_base_plus_offset/sum_rename_ack
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4727_sample_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4783_update_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Sample/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_word_addrgen/root_register_req
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Update/word_access_complete/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Update/word_access_complete/word_0/cr
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Update/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_base_plus_offset/sum_rename_req
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Update/word_access_complete/word_0/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4822_update_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Sample/word_access_start/word_0/rr
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Sample/word_access_start/word_0/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Sample/word_access_start/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Update/word_access_complete/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_word_addrgen/root_register_ack
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_word_addrgen/$exit
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_word_addrgen/root_register_req
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_word_addrgen/$exit
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_word_addrgen/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Update/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_Sample/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_root_address_calculated
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_word_address_calculated
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_update_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Update/word_access_complete/word_0/cr
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/type_cast_4822_Update/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_depth_high_4755_sample_start_
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Sample/word_access_start/word_0/rr
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Sample/word_access_start/word_0/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Update/word_access_complete/word_0/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Update/word_access_complete/word_0/cr
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_base_plus_offset/$exit
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4767_Sample/word_access_start/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/ptr_deref_4779_Update/word_access_complete/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Update/word_access_complete/word_0/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Update/word_access_complete/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Update/$entry
      -- CP-element group 1185: 	 branch_block_stmt_714/assign_stmt_4728_to_assign_stmt_4864/LOAD_pad_4752_Sample/word_access_start/word_0/rr
      -- CP-element group 1185: 	 branch_block_stmt_714/merge_stmt_4711_PhiAck/$exit
      -- 
    cr_9974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => type_cast_4737_inst_req_1); -- 
    cr_10154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => type_cast_4783_inst_req_1); -- 
    rr_9969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => type_cast_4737_inst_req_0); -- 
    rr_10124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => ptr_deref_4779_load_0_req_0); -- 
    cr_9960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => type_cast_4727_inst_req_1); -- 
    rr_9955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => type_cast_4727_inst_req_0); -- 
    cr_10168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => type_cast_4822_inst_req_1); -- 
    cr_10035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => LOAD_depth_high_4755_load_0_req_1); -- 
    cr_10085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => ptr_deref_4767_load_0_req_1); -- 
    rr_10024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => LOAD_depth_high_4755_load_0_req_0); -- 
    cr_10135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => ptr_deref_4779_load_0_req_1); -- 
    rr_10074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => ptr_deref_4767_load_0_req_0); -- 
    cr_10002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => LOAD_pad_4752_load_0_req_1); -- 
    rr_9991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => LOAD_pad_4752_load_0_req_0); -- 
    zeropad3D_cp_element_group_1185: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1185"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1182) & zeropad3D_CP_2152_elements(1183) & zeropad3D_CP_2152_elements(1184);
      gj_zeropad3D_cp_element_group_1185 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1186:  transition  input  bypass 
    -- CP-element group 1186: predecessors 
    -- CP-element group 1186: 	8 
    -- CP-element group 1186: successors 
    -- CP-element group 1186: 	1188 
    -- CP-element group 1186:  members (2) 
      -- CP-element group 1186: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4879/SplitProtocol/Sample/$exit
      -- CP-element group 1186: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4879/SplitProtocol/Sample/ra
      -- 
    ra_13962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4879_inst_ack_0, ack => zeropad3D_CP_2152_elements(1186)); -- 
    -- CP-element group 1187:  transition  input  bypass 
    -- CP-element group 1187: predecessors 
    -- CP-element group 1187: 	8 
    -- CP-element group 1187: successors 
    -- CP-element group 1187: 	1188 
    -- CP-element group 1187:  members (2) 
      -- CP-element group 1187: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4879/SplitProtocol/Update/$exit
      -- CP-element group 1187: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4879/SplitProtocol/Update/ca
      -- 
    ca_13967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4879_inst_ack_1, ack => zeropad3D_CP_2152_elements(1187)); -- 
    -- CP-element group 1188:  join  transition  output  bypass 
    -- CP-element group 1188: predecessors 
    -- CP-element group 1188: 	1186 
    -- CP-element group 1188: 	1187 
    -- CP-element group 1188: successors 
    -- CP-element group 1188: 	1195 
    -- CP-element group 1188:  members (5) 
      -- CP-element group 1188: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/$exit
      -- CP-element group 1188: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/$exit
      -- CP-element group 1188: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4879/$exit
      -- CP-element group 1188: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4879/SplitProtocol/$exit
      -- CP-element group 1188: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_req
      -- 
    phi_stmt_4874_req_13968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4874_req_13968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1188), ack => phi_stmt_4874_req_1); -- 
    zeropad3D_cp_element_group_1188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1186) & zeropad3D_CP_2152_elements(1187);
      gj_zeropad3D_cp_element_group_1188 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1189:  transition  input  bypass 
    -- CP-element group 1189: predecessors 
    -- CP-element group 1189: 	8 
    -- CP-element group 1189: successors 
    -- CP-element group 1189: 	1191 
    -- CP-element group 1189:  members (2) 
      -- CP-element group 1189: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4883/SplitProtocol/Sample/$exit
      -- CP-element group 1189: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4883/SplitProtocol/Sample/ra
      -- 
    ra_13985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4883_inst_ack_0, ack => zeropad3D_CP_2152_elements(1189)); -- 
    -- CP-element group 1190:  transition  input  bypass 
    -- CP-element group 1190: predecessors 
    -- CP-element group 1190: 	8 
    -- CP-element group 1190: successors 
    -- CP-element group 1190: 	1191 
    -- CP-element group 1190:  members (2) 
      -- CP-element group 1190: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4883/SplitProtocol/Update/$exit
      -- CP-element group 1190: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4883/SplitProtocol/Update/ca
      -- 
    ca_13990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4883_inst_ack_1, ack => zeropad3D_CP_2152_elements(1190)); -- 
    -- CP-element group 1191:  join  transition  output  bypass 
    -- CP-element group 1191: predecessors 
    -- CP-element group 1191: 	1189 
    -- CP-element group 1191: 	1190 
    -- CP-element group 1191: successors 
    -- CP-element group 1191: 	1195 
    -- CP-element group 1191:  members (5) 
      -- CP-element group 1191: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/$exit
      -- CP-element group 1191: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/$exit
      -- CP-element group 1191: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4883/$exit
      -- CP-element group 1191: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4883/SplitProtocol/$exit
      -- CP-element group 1191: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_req
      -- 
    phi_stmt_4880_req_13991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4880_req_13991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1191), ack => phi_stmt_4880_req_0); -- 
    zeropad3D_cp_element_group_1191: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1191"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1189) & zeropad3D_CP_2152_elements(1190);
      gj_zeropad3D_cp_element_group_1191 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1192:  transition  input  bypass 
    -- CP-element group 1192: predecessors 
    -- CP-element group 1192: 	8 
    -- CP-element group 1192: successors 
    -- CP-element group 1192: 	1194 
    -- CP-element group 1192:  members (2) 
      -- CP-element group 1192: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/type_cast_4873/SplitProtocol/Sample/$exit
      -- CP-element group 1192: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/type_cast_4873/SplitProtocol/Sample/ra
      -- 
    ra_14008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4873_inst_ack_0, ack => zeropad3D_CP_2152_elements(1192)); -- 
    -- CP-element group 1193:  transition  input  bypass 
    -- CP-element group 1193: predecessors 
    -- CP-element group 1193: 	8 
    -- CP-element group 1193: successors 
    -- CP-element group 1193: 	1194 
    -- CP-element group 1193:  members (2) 
      -- CP-element group 1193: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/type_cast_4873/SplitProtocol/Update/$exit
      -- CP-element group 1193: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/type_cast_4873/SplitProtocol/Update/ca
      -- 
    ca_14013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4873_inst_ack_1, ack => zeropad3D_CP_2152_elements(1193)); -- 
    -- CP-element group 1194:  join  transition  output  bypass 
    -- CP-element group 1194: predecessors 
    -- CP-element group 1194: 	1192 
    -- CP-element group 1194: 	1193 
    -- CP-element group 1194: successors 
    -- CP-element group 1194: 	1195 
    -- CP-element group 1194:  members (5) 
      -- CP-element group 1194: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/$exit
      -- CP-element group 1194: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/$exit
      -- CP-element group 1194: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/type_cast_4873/$exit
      -- CP-element group 1194: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/type_cast_4873/SplitProtocol/$exit
      -- CP-element group 1194: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_req
      -- 
    phi_stmt_4867_req_14014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4867_req_14014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1194), ack => phi_stmt_4867_req_1); -- 
    zeropad3D_cp_element_group_1194: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1194"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1192) & zeropad3D_CP_2152_elements(1193);
      gj_zeropad3D_cp_element_group_1194 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1195:  join  transition  bypass 
    -- CP-element group 1195: predecessors 
    -- CP-element group 1195: 	1188 
    -- CP-element group 1195: 	1191 
    -- CP-element group 1195: 	1194 
    -- CP-element group 1195: successors 
    -- CP-element group 1195: 	1204 
    -- CP-element group 1195:  members (1) 
      -- CP-element group 1195: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1195: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1195"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1188) & zeropad3D_CP_2152_elements(1191) & zeropad3D_CP_2152_elements(1194);
      gj_zeropad3D_cp_element_group_1195 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1196:  transition  input  bypass 
    -- CP-element group 1196: predecessors 
    -- CP-element group 1196: 	701 
    -- CP-element group 1196: successors 
    -- CP-element group 1196: 	1198 
    -- CP-element group 1196:  members (2) 
      -- CP-element group 1196: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4877/SplitProtocol/Sample/$exit
      -- CP-element group 1196: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4877/SplitProtocol/Sample/ra
      -- 
    ra_14034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4877_inst_ack_0, ack => zeropad3D_CP_2152_elements(1196)); -- 
    -- CP-element group 1197:  transition  input  bypass 
    -- CP-element group 1197: predecessors 
    -- CP-element group 1197: 	701 
    -- CP-element group 1197: successors 
    -- CP-element group 1197: 	1198 
    -- CP-element group 1197:  members (2) 
      -- CP-element group 1197: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4877/SplitProtocol/Update/ca
      -- CP-element group 1197: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4877/SplitProtocol/Update/$exit
      -- 
    ca_14039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4877_inst_ack_1, ack => zeropad3D_CP_2152_elements(1197)); -- 
    -- CP-element group 1198:  join  transition  output  bypass 
    -- CP-element group 1198: predecessors 
    -- CP-element group 1198: 	1196 
    -- CP-element group 1198: 	1197 
    -- CP-element group 1198: successors 
    -- CP-element group 1198: 	1203 
    -- CP-element group 1198:  members (5) 
      -- CP-element group 1198: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_req
      -- CP-element group 1198: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4877/SplitProtocol/$exit
      -- CP-element group 1198: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/type_cast_4877/$exit
      -- CP-element group 1198: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/$exit
      -- CP-element group 1198: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4874/phi_stmt_4874_sources/$exit
      -- 
    phi_stmt_4874_req_14040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4874_req_14040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1198), ack => phi_stmt_4874_req_0); -- 
    zeropad3D_cp_element_group_1198: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1198"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1196) & zeropad3D_CP_2152_elements(1197);
      gj_zeropad3D_cp_element_group_1198 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1199:  transition  input  bypass 
    -- CP-element group 1199: predecessors 
    -- CP-element group 1199: 	701 
    -- CP-element group 1199: successors 
    -- CP-element group 1199: 	1201 
    -- CP-element group 1199:  members (2) 
      -- CP-element group 1199: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4885/SplitProtocol/Sample/ra
      -- CP-element group 1199: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4885/SplitProtocol/Sample/$exit
      -- 
    ra_14057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4885_inst_ack_0, ack => zeropad3D_CP_2152_elements(1199)); -- 
    -- CP-element group 1200:  transition  input  bypass 
    -- CP-element group 1200: predecessors 
    -- CP-element group 1200: 	701 
    -- CP-element group 1200: successors 
    -- CP-element group 1200: 	1201 
    -- CP-element group 1200:  members (2) 
      -- CP-element group 1200: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4885/SplitProtocol/Update/ca
      -- CP-element group 1200: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4885/SplitProtocol/Update/$exit
      -- 
    ca_14062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4885_inst_ack_1, ack => zeropad3D_CP_2152_elements(1200)); -- 
    -- CP-element group 1201:  join  transition  output  bypass 
    -- CP-element group 1201: predecessors 
    -- CP-element group 1201: 	1199 
    -- CP-element group 1201: 	1200 
    -- CP-element group 1201: successors 
    -- CP-element group 1201: 	1203 
    -- CP-element group 1201:  members (5) 
      -- CP-element group 1201: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_req
      -- CP-element group 1201: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4885/SplitProtocol/$exit
      -- CP-element group 1201: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/type_cast_4885/$exit
      -- CP-element group 1201: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/phi_stmt_4880_sources/$exit
      -- CP-element group 1201: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4880/$exit
      -- 
    phi_stmt_4880_req_14063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4880_req_14063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1201), ack => phi_stmt_4880_req_1); -- 
    zeropad3D_cp_element_group_1201: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1201"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1199) & zeropad3D_CP_2152_elements(1200);
      gj_zeropad3D_cp_element_group_1201 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1202:  transition  output  delay-element  bypass 
    -- CP-element group 1202: predecessors 
    -- CP-element group 1202: 	701 
    -- CP-element group 1202: successors 
    -- CP-element group 1202: 	1203 
    -- CP-element group 1202:  members (4) 
      -- CP-element group 1202: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/$exit
      -- CP-element group 1202: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4867/$exit
      -- CP-element group 1202: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_req
      -- CP-element group 1202: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4867/phi_stmt_4867_sources/type_cast_4871_konst_delay_trans
      -- 
    phi_stmt_4867_req_14071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4867_req_14071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1202), ack => phi_stmt_4867_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(1202) is a control-delay.
    cp_element_1202_delay: control_delay_element  generic map(name => " 1202_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(701), ack => zeropad3D_CP_2152_elements(1202), clk => clk, reset =>reset);
    -- CP-element group 1203:  join  transition  bypass 
    -- CP-element group 1203: predecessors 
    -- CP-element group 1203: 	1198 
    -- CP-element group 1203: 	1201 
    -- CP-element group 1203: 	1202 
    -- CP-element group 1203: successors 
    -- CP-element group 1203: 	1204 
    -- CP-element group 1203:  members (1) 
      -- CP-element group 1203: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1203: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1203"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1198) & zeropad3D_CP_2152_elements(1201) & zeropad3D_CP_2152_elements(1202);
      gj_zeropad3D_cp_element_group_1203 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1204:  merge  fork  transition  place  bypass 
    -- CP-element group 1204: predecessors 
    -- CP-element group 1204: 	1195 
    -- CP-element group 1204: 	1203 
    -- CP-element group 1204: successors 
    -- CP-element group 1204: 	1205 
    -- CP-element group 1204: 	1206 
    -- CP-element group 1204: 	1207 
    -- CP-element group 1204:  members (2) 
      -- CP-element group 1204: 	 branch_block_stmt_714/merge_stmt_4866_PhiReqMerge
      -- CP-element group 1204: 	 branch_block_stmt_714/merge_stmt_4866_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1204) <= OrReduce(zeropad3D_CP_2152_elements(1195) & zeropad3D_CP_2152_elements(1203));
    -- CP-element group 1205:  transition  input  bypass 
    -- CP-element group 1205: predecessors 
    -- CP-element group 1205: 	1204 
    -- CP-element group 1205: successors 
    -- CP-element group 1205: 	1208 
    -- CP-element group 1205:  members (1) 
      -- CP-element group 1205: 	 branch_block_stmt_714/merge_stmt_4866_PhiAck/phi_stmt_4867_ack
      -- 
    phi_stmt_4867_ack_14076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4867_ack_0, ack => zeropad3D_CP_2152_elements(1205)); -- 
    -- CP-element group 1206:  transition  input  bypass 
    -- CP-element group 1206: predecessors 
    -- CP-element group 1206: 	1204 
    -- CP-element group 1206: successors 
    -- CP-element group 1206: 	1208 
    -- CP-element group 1206:  members (1) 
      -- CP-element group 1206: 	 branch_block_stmt_714/merge_stmt_4866_PhiAck/phi_stmt_4874_ack
      -- 
    phi_stmt_4874_ack_14077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4874_ack_0, ack => zeropad3D_CP_2152_elements(1206)); -- 
    -- CP-element group 1207:  transition  input  bypass 
    -- CP-element group 1207: predecessors 
    -- CP-element group 1207: 	1204 
    -- CP-element group 1207: successors 
    -- CP-element group 1207: 	1208 
    -- CP-element group 1207:  members (1) 
      -- CP-element group 1207: 	 branch_block_stmt_714/merge_stmt_4866_PhiAck/phi_stmt_4880_ack
      -- 
    phi_stmt_4880_ack_14078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4880_ack_0, ack => zeropad3D_CP_2152_elements(1207)); -- 
    -- CP-element group 1208:  join  fork  transition  place  output  bypass 
    -- CP-element group 1208: predecessors 
    -- CP-element group 1208: 	1205 
    -- CP-element group 1208: 	1206 
    -- CP-element group 1208: 	1207 
    -- CP-element group 1208: successors 
    -- CP-element group 1208: 	702 
    -- CP-element group 1208: 	703 
    -- CP-element group 1208:  members (10) 
      -- CP-element group 1208: 	 branch_block_stmt_714/merge_stmt_4866__exit__
      -- CP-element group 1208: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898__entry__
      -- CP-element group 1208: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/type_cast_4890_Update/$entry
      -- CP-element group 1208: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/type_cast_4890_sample_start_
      -- CP-element group 1208: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/type_cast_4890_Update/cr
      -- CP-element group 1208: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/$entry
      -- CP-element group 1208: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/type_cast_4890_Sample/rr
      -- CP-element group 1208: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/type_cast_4890_Sample/$entry
      -- CP-element group 1208: 	 branch_block_stmt_714/assign_stmt_4891_to_assign_stmt_4898/type_cast_4890_update_start_
      -- CP-element group 1208: 	 branch_block_stmt_714/merge_stmt_4866_PhiAck/$exit
      -- 
    cr_10185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1208), ack => type_cast_4890_inst_req_1); -- 
    rr_10180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1208), ack => type_cast_4890_inst_req_0); -- 
    zeropad3D_cp_element_group_1208: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1208"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1205) & zeropad3D_CP_2152_elements(1206) & zeropad3D_CP_2152_elements(1207);
      gj_zeropad3D_cp_element_group_1208 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1209:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1209: predecessors 
    -- CP-element group 1209: 	704 
    -- CP-element group 1209: 	711 
    -- CP-element group 1209: 	714 
    -- CP-element group 1209: 	721 
    -- CP-element group 1209: successors 
    -- CP-element group 1209: 	722 
    -- CP-element group 1209: 	723 
    -- CP-element group 1209: 	724 
    -- CP-element group 1209: 	725 
    -- CP-element group 1209: 	728 
    -- CP-element group 1209: 	730 
    -- CP-element group 1209: 	732 
    -- CP-element group 1209: 	734 
    -- CP-element group 1209:  members (33) 
      -- CP-element group 1209: 	 branch_block_stmt_714/merge_stmt_4976__exit__
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032__entry__
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/$entry
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4980_sample_start_
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4980_update_start_
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4980_Sample/$entry
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4980_Sample/rr
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4980_Update/$entry
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4980_Update/cr
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4985_sample_start_
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4985_update_start_
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4985_Sample/$entry
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4985_Sample/rr
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4985_Update/$entry
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_4985_Update/cr
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_5019_update_start_
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_5019_Update/$entry
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/type_cast_5019_Update/cr
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/addr_of_5026_update_start_
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_final_index_sum_regn_update_start
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_final_index_sum_regn_Update/$entry
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/array_obj_ref_5025_final_index_sum_regn_Update/req
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/addr_of_5026_complete/$entry
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/addr_of_5026_complete/req
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_update_start_
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Update/$entry
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Update/word_access_complete/$entry
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Update/word_access_complete/word_0/$entry
      -- CP-element group 1209: 	 branch_block_stmt_714/assign_stmt_4981_to_assign_stmt_5032/ptr_deref_5029_Update/word_access_complete/word_0/cr
      -- CP-element group 1209: 	 branch_block_stmt_714/merge_stmt_4976_PhiReqMerge
      -- CP-element group 1209: 	 branch_block_stmt_714/merge_stmt_4976_PhiAck/dummy
      -- CP-element group 1209: 	 branch_block_stmt_714/merge_stmt_4976_PhiAck/$exit
      -- CP-element group 1209: 	 branch_block_stmt_714/merge_stmt_4976_PhiAck/$entry
      -- 
    rr_10390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1209), ack => type_cast_4980_inst_req_0); -- 
    cr_10395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1209), ack => type_cast_4980_inst_req_1); -- 
    rr_10404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1209), ack => type_cast_4985_inst_req_0); -- 
    cr_10409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1209), ack => type_cast_4985_inst_req_1); -- 
    cr_10423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1209), ack => type_cast_5019_inst_req_1); -- 
    req_10454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1209), ack => array_obj_ref_5025_index_offset_req_1); -- 
    req_10469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1209), ack => addr_of_5026_final_reg_req_1); -- 
    cr_10519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1209), ack => ptr_deref_5029_store_0_req_1); -- 
    zeropad3D_CP_2152_elements(1209) <= OrReduce(zeropad3D_CP_2152_elements(704) & zeropad3D_CP_2152_elements(711) & zeropad3D_CP_2152_elements(714) & zeropad3D_CP_2152_elements(721));
    -- CP-element group 1210:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1210: predecessors 
    -- CP-element group 1210: 	735 
    -- CP-element group 1210: 	755 
    -- CP-element group 1210: successors 
    -- CP-element group 1210: 	756 
    -- CP-element group 1210: 	757 
    -- CP-element group 1210:  members (13) 
      -- CP-element group 1210: 	 branch_block_stmt_714/merge_stmt_5141__exit__
      -- CP-element group 1210: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159__entry__
      -- CP-element group 1210: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/$entry
      -- CP-element group 1210: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/type_cast_5145_sample_start_
      -- CP-element group 1210: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/type_cast_5145_update_start_
      -- CP-element group 1210: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/type_cast_5145_Sample/$entry
      -- CP-element group 1210: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/type_cast_5145_Sample/rr
      -- CP-element group 1210: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/type_cast_5145_Update/$entry
      -- CP-element group 1210: 	 branch_block_stmt_714/assign_stmt_5146_to_assign_stmt_5159/type_cast_5145_Update/cr
      -- CP-element group 1210: 	 branch_block_stmt_714/merge_stmt_5141_PhiAck/dummy
      -- CP-element group 1210: 	 branch_block_stmt_714/merge_stmt_5141_PhiAck/$exit
      -- CP-element group 1210: 	 branch_block_stmt_714/merge_stmt_5141_PhiAck/$entry
      -- CP-element group 1210: 	 branch_block_stmt_714/merge_stmt_5141_PhiReqMerge
      -- 
    rr_10768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1210), ack => type_cast_5145_inst_req_0); -- 
    cr_10773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1210), ack => type_cast_5145_inst_req_1); -- 
    zeropad3D_CP_2152_elements(1210) <= OrReduce(zeropad3D_CP_2152_elements(735) & zeropad3D_CP_2152_elements(755));
    -- CP-element group 1211:  transition  output  delay-element  bypass 
    -- CP-element group 1211: predecessors 
    -- CP-element group 1211: 	777 
    -- CP-element group 1211: successors 
    -- CP-element group 1211: 	1218 
    -- CP-element group 1211:  members (4) 
      -- CP-element group 1211: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5247/$exit
      -- CP-element group 1211: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_req
      -- CP-element group 1211: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/type_cast_5253_konst_delay_trans
      -- CP-element group 1211: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/$exit
      -- 
    phi_stmt_5247_req_14189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_5247_req_14189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1211), ack => phi_stmt_5247_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(1211) is a control-delay.
    cp_element_1211_delay: control_delay_element  generic map(name => " 1211_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(777), ack => zeropad3D_CP_2152_elements(1211), clk => clk, reset =>reset);
    -- CP-element group 1212:  transition  input  bypass 
    -- CP-element group 1212: predecessors 
    -- CP-element group 1212: 	777 
    -- CP-element group 1212: successors 
    -- CP-element group 1212: 	1214 
    -- CP-element group 1212:  members (2) 
      -- CP-element group 1212: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5259/SplitProtocol/Sample/ra
      -- CP-element group 1212: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5259/SplitProtocol/Sample/$exit
      -- 
    ra_14206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5259_inst_ack_0, ack => zeropad3D_CP_2152_elements(1212)); -- 
    -- CP-element group 1213:  transition  input  bypass 
    -- CP-element group 1213: predecessors 
    -- CP-element group 1213: 	777 
    -- CP-element group 1213: successors 
    -- CP-element group 1213: 	1214 
    -- CP-element group 1213:  members (2) 
      -- CP-element group 1213: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5259/SplitProtocol/Update/ca
      -- CP-element group 1213: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5259/SplitProtocol/Update/$exit
      -- 
    ca_14211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5259_inst_ack_1, ack => zeropad3D_CP_2152_elements(1213)); -- 
    -- CP-element group 1214:  join  transition  output  bypass 
    -- CP-element group 1214: predecessors 
    -- CP-element group 1214: 	1212 
    -- CP-element group 1214: 	1213 
    -- CP-element group 1214: successors 
    -- CP-element group 1214: 	1218 
    -- CP-element group 1214:  members (5) 
      -- CP-element group 1214: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_req
      -- CP-element group 1214: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5259/SplitProtocol/$exit
      -- CP-element group 1214: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5259/$exit
      -- CP-element group 1214: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/$exit
      -- CP-element group 1214: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5254/$exit
      -- 
    phi_stmt_5254_req_14212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_5254_req_14212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1214), ack => phi_stmt_5254_req_1); -- 
    zeropad3D_cp_element_group_1214: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1214"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1212) & zeropad3D_CP_2152_elements(1213);
      gj_zeropad3D_cp_element_group_1214 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1215:  transition  input  bypass 
    -- CP-element group 1215: predecessors 
    -- CP-element group 1215: 	777 
    -- CP-element group 1215: successors 
    -- CP-element group 1215: 	1217 
    -- CP-element group 1215:  members (2) 
      -- CP-element group 1215: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5263/SplitProtocol/Sample/$exit
      -- CP-element group 1215: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5263/SplitProtocol/Sample/ra
      -- 
    ra_14229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5263_inst_ack_0, ack => zeropad3D_CP_2152_elements(1215)); -- 
    -- CP-element group 1216:  transition  input  bypass 
    -- CP-element group 1216: predecessors 
    -- CP-element group 1216: 	777 
    -- CP-element group 1216: successors 
    -- CP-element group 1216: 	1217 
    -- CP-element group 1216:  members (2) 
      -- CP-element group 1216: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5263/SplitProtocol/Update/$exit
      -- CP-element group 1216: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5263/SplitProtocol/Update/ca
      -- 
    ca_14234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5263_inst_ack_1, ack => zeropad3D_CP_2152_elements(1216)); -- 
    -- CP-element group 1217:  join  transition  output  bypass 
    -- CP-element group 1217: predecessors 
    -- CP-element group 1217: 	1215 
    -- CP-element group 1217: 	1216 
    -- CP-element group 1217: successors 
    -- CP-element group 1217: 	1218 
    -- CP-element group 1217:  members (5) 
      -- CP-element group 1217: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5263/SplitProtocol/$exit
      -- CP-element group 1217: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5263/$exit
      -- CP-element group 1217: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/$exit
      -- CP-element group 1217: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/$exit
      -- CP-element group 1217: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_req
      -- 
    phi_stmt_5260_req_14235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_5260_req_14235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1217), ack => phi_stmt_5260_req_0); -- 
    zeropad3D_cp_element_group_1217: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1217"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1215) & zeropad3D_CP_2152_elements(1216);
      gj_zeropad3D_cp_element_group_1217 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1218:  join  transition  bypass 
    -- CP-element group 1218: predecessors 
    -- CP-element group 1218: 	1211 
    -- CP-element group 1218: 	1214 
    -- CP-element group 1218: 	1217 
    -- CP-element group 1218: successors 
    -- CP-element group 1218: 	1229 
    -- CP-element group 1218:  members (1) 
      -- CP-element group 1218: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1218: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1218"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1211) & zeropad3D_CP_2152_elements(1214) & zeropad3D_CP_2152_elements(1217);
      gj_zeropad3D_cp_element_group_1218 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1219:  transition  input  bypass 
    -- CP-element group 1219: predecessors 
    -- CP-element group 1219: 	758 
    -- CP-element group 1219: successors 
    -- CP-element group 1219: 	1221 
    -- CP-element group 1219:  members (2) 
      -- CP-element group 1219: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/type_cast_5250/SplitProtocol/Sample/ra
      -- CP-element group 1219: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/type_cast_5250/SplitProtocol/Sample/$exit
      -- 
    ra_14255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5250_inst_ack_0, ack => zeropad3D_CP_2152_elements(1219)); -- 
    -- CP-element group 1220:  transition  input  bypass 
    -- CP-element group 1220: predecessors 
    -- CP-element group 1220: 	758 
    -- CP-element group 1220: successors 
    -- CP-element group 1220: 	1221 
    -- CP-element group 1220:  members (2) 
      -- CP-element group 1220: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/type_cast_5250/SplitProtocol/Update/ca
      -- CP-element group 1220: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/type_cast_5250/SplitProtocol/Update/$exit
      -- 
    ca_14260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5250_inst_ack_1, ack => zeropad3D_CP_2152_elements(1220)); -- 
    -- CP-element group 1221:  join  transition  output  bypass 
    -- CP-element group 1221: predecessors 
    -- CP-element group 1221: 	1219 
    -- CP-element group 1221: 	1220 
    -- CP-element group 1221: successors 
    -- CP-element group 1221: 	1228 
    -- CP-element group 1221:  members (5) 
      -- CP-element group 1221: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/type_cast_5250/$exit
      -- CP-element group 1221: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/$exit
      -- CP-element group 1221: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/$exit
      -- CP-element group 1221: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_req
      -- CP-element group 1221: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5247/phi_stmt_5247_sources/type_cast_5250/SplitProtocol/$exit
      -- 
    phi_stmt_5247_req_14261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_5247_req_14261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1221), ack => phi_stmt_5247_req_0); -- 
    zeropad3D_cp_element_group_1221: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1221"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1219) & zeropad3D_CP_2152_elements(1220);
      gj_zeropad3D_cp_element_group_1221 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1222:  transition  input  bypass 
    -- CP-element group 1222: predecessors 
    -- CP-element group 1222: 	758 
    -- CP-element group 1222: successors 
    -- CP-element group 1222: 	1224 
    -- CP-element group 1222:  members (2) 
      -- CP-element group 1222: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5257/SplitProtocol/Sample/ra
      -- CP-element group 1222: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5257/SplitProtocol/Sample/$exit
      -- 
    ra_14278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5257_inst_ack_0, ack => zeropad3D_CP_2152_elements(1222)); -- 
    -- CP-element group 1223:  transition  input  bypass 
    -- CP-element group 1223: predecessors 
    -- CP-element group 1223: 	758 
    -- CP-element group 1223: successors 
    -- CP-element group 1223: 	1224 
    -- CP-element group 1223:  members (2) 
      -- CP-element group 1223: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5257/SplitProtocol/Update/ca
      -- CP-element group 1223: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5257/SplitProtocol/Update/$exit
      -- 
    ca_14283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5257_inst_ack_1, ack => zeropad3D_CP_2152_elements(1223)); -- 
    -- CP-element group 1224:  join  transition  output  bypass 
    -- CP-element group 1224: predecessors 
    -- CP-element group 1224: 	1222 
    -- CP-element group 1224: 	1223 
    -- CP-element group 1224: successors 
    -- CP-element group 1224: 	1228 
    -- CP-element group 1224:  members (5) 
      -- CP-element group 1224: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_req
      -- CP-element group 1224: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5257/SplitProtocol/$exit
      -- CP-element group 1224: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/type_cast_5257/$exit
      -- CP-element group 1224: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/phi_stmt_5254_sources/$exit
      -- CP-element group 1224: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5254/$exit
      -- 
    phi_stmt_5254_req_14284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_5254_req_14284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1224), ack => phi_stmt_5254_req_0); -- 
    zeropad3D_cp_element_group_1224: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1224"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1222) & zeropad3D_CP_2152_elements(1223);
      gj_zeropad3D_cp_element_group_1224 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1224), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1225:  transition  input  bypass 
    -- CP-element group 1225: predecessors 
    -- CP-element group 1225: 	758 
    -- CP-element group 1225: successors 
    -- CP-element group 1225: 	1227 
    -- CP-element group 1225:  members (2) 
      -- CP-element group 1225: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5265/SplitProtocol/Sample/$exit
      -- CP-element group 1225: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5265/SplitProtocol/Sample/ra
      -- 
    ra_14301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5265_inst_ack_0, ack => zeropad3D_CP_2152_elements(1225)); -- 
    -- CP-element group 1226:  transition  input  bypass 
    -- CP-element group 1226: predecessors 
    -- CP-element group 1226: 	758 
    -- CP-element group 1226: successors 
    -- CP-element group 1226: 	1227 
    -- CP-element group 1226:  members (2) 
      -- CP-element group 1226: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5265/SplitProtocol/Update/ca
      -- CP-element group 1226: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5265/SplitProtocol/Update/$exit
      -- 
    ca_14306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5265_inst_ack_1, ack => zeropad3D_CP_2152_elements(1226)); -- 
    -- CP-element group 1227:  join  transition  output  bypass 
    -- CP-element group 1227: predecessors 
    -- CP-element group 1227: 	1225 
    -- CP-element group 1227: 	1226 
    -- CP-element group 1227: successors 
    -- CP-element group 1227: 	1228 
    -- CP-element group 1227:  members (5) 
      -- CP-element group 1227: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5265/$exit
      -- CP-element group 1227: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/type_cast_5265/SplitProtocol/$exit
      -- CP-element group 1227: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_sources/$exit
      -- CP-element group 1227: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/$exit
      -- CP-element group 1227: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5260/phi_stmt_5260_req
      -- 
    phi_stmt_5260_req_14307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_5260_req_14307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1227), ack => phi_stmt_5260_req_1); -- 
    zeropad3D_cp_element_group_1227: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1227"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1225) & zeropad3D_CP_2152_elements(1226);
      gj_zeropad3D_cp_element_group_1227 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1228:  join  transition  bypass 
    -- CP-element group 1228: predecessors 
    -- CP-element group 1228: 	1221 
    -- CP-element group 1228: 	1224 
    -- CP-element group 1228: 	1227 
    -- CP-element group 1228: successors 
    -- CP-element group 1228: 	1229 
    -- CP-element group 1228:  members (1) 
      -- CP-element group 1228: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1228: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1228"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1221) & zeropad3D_CP_2152_elements(1224) & zeropad3D_CP_2152_elements(1227);
      gj_zeropad3D_cp_element_group_1228 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1229:  merge  fork  transition  place  bypass 
    -- CP-element group 1229: predecessors 
    -- CP-element group 1229: 	1218 
    -- CP-element group 1229: 	1228 
    -- CP-element group 1229: successors 
    -- CP-element group 1229: 	1230 
    -- CP-element group 1229: 	1231 
    -- CP-element group 1229: 	1232 
    -- CP-element group 1229:  members (2) 
      -- CP-element group 1229: 	 branch_block_stmt_714/merge_stmt_5246_PhiAck/$entry
      -- CP-element group 1229: 	 branch_block_stmt_714/merge_stmt_5246_PhiReqMerge
      -- 
    zeropad3D_CP_2152_elements(1229) <= OrReduce(zeropad3D_CP_2152_elements(1218) & zeropad3D_CP_2152_elements(1228));
    -- CP-element group 1230:  transition  input  bypass 
    -- CP-element group 1230: predecessors 
    -- CP-element group 1230: 	1229 
    -- CP-element group 1230: successors 
    -- CP-element group 1230: 	1233 
    -- CP-element group 1230:  members (1) 
      -- CP-element group 1230: 	 branch_block_stmt_714/merge_stmt_5246_PhiAck/phi_stmt_5247_ack
      -- 
    phi_stmt_5247_ack_14312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_5247_ack_0, ack => zeropad3D_CP_2152_elements(1230)); -- 
    -- CP-element group 1231:  transition  input  bypass 
    -- CP-element group 1231: predecessors 
    -- CP-element group 1231: 	1229 
    -- CP-element group 1231: successors 
    -- CP-element group 1231: 	1233 
    -- CP-element group 1231:  members (1) 
      -- CP-element group 1231: 	 branch_block_stmt_714/merge_stmt_5246_PhiAck/phi_stmt_5254_ack
      -- 
    phi_stmt_5254_ack_14313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_5254_ack_0, ack => zeropad3D_CP_2152_elements(1231)); -- 
    -- CP-element group 1232:  transition  input  bypass 
    -- CP-element group 1232: predecessors 
    -- CP-element group 1232: 	1229 
    -- CP-element group 1232: successors 
    -- CP-element group 1232: 	1233 
    -- CP-element group 1232:  members (1) 
      -- CP-element group 1232: 	 branch_block_stmt_714/merge_stmt_5246_PhiAck/phi_stmt_5260_ack
      -- 
    phi_stmt_5260_ack_14314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_5260_ack_0, ack => zeropad3D_CP_2152_elements(1232)); -- 
    -- CP-element group 1233:  join  transition  bypass 
    -- CP-element group 1233: predecessors 
    -- CP-element group 1233: 	1230 
    -- CP-element group 1233: 	1231 
    -- CP-element group 1233: 	1232 
    -- CP-element group 1233: successors 
    -- CP-element group 1233: 	8 
    -- CP-element group 1233:  members (1) 
      -- CP-element group 1233: 	 branch_block_stmt_714/merge_stmt_5246_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1233: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1233"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1230) & zeropad3D_CP_2152_elements(1231) & zeropad3D_CP_2152_elements(1232);
      gj_zeropad3D_cp_element_group_1233 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1233), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1059_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1143_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1168_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1394_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1409_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1433_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1459_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1617_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1700_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1725_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1944_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1959_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1983_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2009_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2173_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2256_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2281_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2521_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2536_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2560_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2586_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2743_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2826_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2851_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3070_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3085_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3109_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3135_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3305_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3388_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3413_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3659_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3674_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3698_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3724_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3887_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3970_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3995_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4226_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4241_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4265_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4291_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4449_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4532_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4557_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4797_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4812_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4836_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4862_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_5013_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_5096_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_5121_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_829_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_844_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_868_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_894_wire : std_logic_vector(31 downto 0);
    signal LOAD_col_high_1234_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_1234_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_1556_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_1556_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_1791_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_1791_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_2106_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_2106_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_2347_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_2347_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_2682_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_2682_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_2917_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_2917_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_3238_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_3238_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_3479_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_3479_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_3826_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_3826_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4061_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4061_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4382_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4382_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4623_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4623_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4952_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4952_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_5187_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_5187_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_782_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_782_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_992_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_992_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_1352_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_1352_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_1902_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_1902_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_2479_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_2479_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_3028_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_3028_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_3617_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_3617_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_4184_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_4184_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_4755_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_4755_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_779_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_779_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_1349_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_1349_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_1899_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_1899_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_2476_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_2476_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_3025_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_3025_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_3614_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_3614_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_4181_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_4181_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_4752_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_4752_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_776_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_776_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_1278_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_1278_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_1505_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_1505_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_1828_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_1828_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_2055_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_2055_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_2391_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_2391_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_2631_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_2631_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_2954_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_2954_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_3181_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_3181_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_3523_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_3523_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_3769_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_3769_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_4098_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_4098_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_4337_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_4337_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_4667_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_4667_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_4907_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_4907_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_5224_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_5224_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_941_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_941_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom1002_3424_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1002_3424_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1177_3898_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1177_3898_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1220_3981_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1220_3981_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1225_4006_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1225_4006_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom130_1154_resized : std_logic_vector(13 downto 0);
    signal R_idxprom130_1154_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom135_1179_resized : std_logic_vector(13 downto 0);
    signal R_idxprom135_1179_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1395_4460_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1395_4460_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1438_4543_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1438_4543_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1443_4568_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1443_4568_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1615_5024_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1615_5024_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1658_5107_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1658_5107_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1663_5132_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1663_5132_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom298_1628_resized : std_logic_vector(13 downto 0);
    signal R_idxprom298_1628_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom341_1711_resized : std_logic_vector(13 downto 0);
    signal R_idxprom341_1711_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom346_1736_resized : std_logic_vector(13 downto 0);
    signal R_idxprom346_1736_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom515_2184_resized : std_logic_vector(13 downto 0);
    signal R_idxprom515_2184_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom558_2267_resized : std_logic_vector(13 downto 0);
    signal R_idxprom558_2267_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom563_2292_resized : std_logic_vector(13 downto 0);
    signal R_idxprom563_2292_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom736_2754_resized : std_logic_vector(13 downto 0);
    signal R_idxprom736_2754_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom779_2837_resized : std_logic_vector(13 downto 0);
    signal R_idxprom779_2837_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom784_2862_resized : std_logic_vector(13 downto 0);
    signal R_idxprom784_2862_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom954_3316_resized : std_logic_vector(13 downto 0);
    signal R_idxprom954_3316_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom997_3399_resized : std_logic_vector(13 downto 0);
    signal R_idxprom997_3399_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1071_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1071_scaled : std_logic_vector(13 downto 0);
    signal STORE_col_high_752_data_0 : std_logic_vector(7 downto 0);
    signal STORE_col_high_752_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_depth_high_771_data_0 : std_logic_vector(7 downto 0);
    signal STORE_depth_high_771_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_row_high_733_data_0 : std_logic_vector(7 downto 0);
    signal STORE_row_high_733_word_address_0 : std_logic_vector(0 downto 0);
    signal add1009_3444 : std_logic_vector(31 downto 0);
    signal add1017_3464 : std_logic_vector(15 downto 0);
    signal add102_1111 : std_logic_vector(31 downto 0);
    signal add1030_3495 : std_logic_vector(31 downto 0);
    signal add1047_3545 : std_logic_vector(31 downto 0);
    signal add111_1116 : std_logic_vector(31 downto 0);
    signal add1138_3791 : std_logic_vector(31 downto 0);
    signal add1155_3836 : std_logic_vector(31 downto 0);
    signal add1168_3875 : std_logic_vector(31 downto 0);
    signal add1174_3880 : std_logic_vector(31 downto 0);
    signal add1192_3938 : std_logic_vector(31 downto 0);
    signal add1201_3943 : std_logic_vector(31 downto 0);
    signal add1211_3958 : std_logic_vector(31 downto 0);
    signal add1217_3963 : std_logic_vector(31 downto 0);
    signal add121_1131 : std_logic_vector(31 downto 0);
    signal add1232_4026 : std_logic_vector(31 downto 0);
    signal add1240_4046 : std_logic_vector(15 downto 0);
    signal add1252_4071 : std_logic_vector(31 downto 0);
    signal add1269_4120 : std_logic_vector(31 downto 0);
    signal add127_1136 : std_logic_vector(31 downto 0);
    signal add1355_4347 : std_logic_vector(31 downto 0);
    signal add1373_4398 : std_logic_vector(31 downto 0);
    signal add1386_4437 : std_logic_vector(31 downto 0);
    signal add1392_4442 : std_logic_vector(31 downto 0);
    signal add140_1199 : std_logic_vector(31 downto 0);
    signal add1410_4500 : std_logic_vector(31 downto 0);
    signal add1419_4505 : std_logic_vector(31 downto 0);
    signal add1429_4520 : std_logic_vector(31 downto 0);
    signal add1435_4525 : std_logic_vector(31 downto 0);
    signal add1450_4588 : std_logic_vector(31 downto 0);
    signal add1458_4608 : std_logic_vector(15 downto 0);
    signal add1471_4639 : std_logic_vector(31 downto 0);
    signal add1486_4677 : std_logic_vector(31 downto 0);
    signal add148_1219 : std_logic_vector(15 downto 0);
    signal add1576_4917 : std_logic_vector(31 downto 0);
    signal add1593_4962 : std_logic_vector(31 downto 0);
    signal add159_1250 : std_logic_vector(31 downto 0);
    signal add1606_5001 : std_logic_vector(31 downto 0);
    signal add1612_5006 : std_logic_vector(31 downto 0);
    signal add1630_5064 : std_logic_vector(31 downto 0);
    signal add1639_5069 : std_logic_vector(31 downto 0);
    signal add1649_5084 : std_logic_vector(31 downto 0);
    signal add1655_5089 : std_logic_vector(31 downto 0);
    signal add1670_5152 : std_logic_vector(31 downto 0);
    signal add1678_5172 : std_logic_vector(15 downto 0);
    signal add1690_5197 : std_logic_vector(31 downto 0);
    signal add1705_5234 : std_logic_vector(31 downto 0);
    signal add175_1294 : std_logic_vector(31 downto 0);
    signal add259_1521 : std_logic_vector(31 downto 0);
    signal add276_1566 : std_logic_vector(31 downto 0);
    signal add289_1605 : std_logic_vector(31 downto 0);
    signal add295_1610 : std_logic_vector(31 downto 0);
    signal add313_1668 : std_logic_vector(31 downto 0);
    signal add322_1673 : std_logic_vector(31 downto 0);
    signal add332_1688 : std_logic_vector(31 downto 0);
    signal add338_1693 : std_logic_vector(31 downto 0);
    signal add353_1756 : std_logic_vector(31 downto 0);
    signal add361_1776 : std_logic_vector(15 downto 0);
    signal add373_1801 : std_logic_vector(31 downto 0);
    signal add389_1844 : std_logic_vector(31 downto 0);
    signal add475_2071 : std_logic_vector(31 downto 0);
    signal add493_2122 : std_logic_vector(31 downto 0);
    signal add506_2161 : std_logic_vector(31 downto 0);
    signal add512_2166 : std_logic_vector(31 downto 0);
    signal add530_2224 : std_logic_vector(31 downto 0);
    signal add539_2229 : std_logic_vector(31 downto 0);
    signal add549_2244 : std_logic_vector(31 downto 0);
    signal add555_2249 : std_logic_vector(31 downto 0);
    signal add570_2312 : std_logic_vector(31 downto 0);
    signal add578_2332 : std_logic_vector(15 downto 0);
    signal add591_2363 : std_logic_vector(31 downto 0);
    signal add607_2407 : std_logic_vector(31 downto 0);
    signal add697_2647 : std_logic_vector(31 downto 0);
    signal add714_2692 : std_logic_vector(31 downto 0);
    signal add727_2731 : std_logic_vector(31 downto 0);
    signal add733_2736 : std_logic_vector(31 downto 0);
    signal add73_1008 : std_logic_vector(31 downto 0);
    signal add751_2794 : std_logic_vector(31 downto 0);
    signal add760_2799 : std_logic_vector(31 downto 0);
    signal add770_2814 : std_logic_vector(31 downto 0);
    signal add776_2819 : std_logic_vector(31 downto 0);
    signal add791_2882 : std_logic_vector(31 downto 0);
    signal add799_2902 : std_logic_vector(15 downto 0);
    signal add811_2927 : std_logic_vector(31 downto 0);
    signal add827_2970 : std_logic_vector(31 downto 0);
    signal add84_1047 : std_logic_vector(31 downto 0);
    signal add90_1052 : std_logic_vector(31 downto 0);
    signal add914_3203 : std_logic_vector(31 downto 0);
    signal add932_3254 : std_logic_vector(31 downto 0);
    signal add945_3293 : std_logic_vector(31 downto 0);
    signal add951_3298 : std_logic_vector(31 downto 0);
    signal add969_3356 : std_logic_vector(31 downto 0);
    signal add978_3361 : std_logic_vector(31 downto 0);
    signal add988_3376 : std_logic_vector(31 downto 0);
    signal add994_3381 : std_logic_vector(31 downto 0);
    signal add_957 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1072_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1180_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1180_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1180_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1180_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1180_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1180_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1629_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1629_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1629_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1629_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1629_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1629_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1712_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1712_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1712_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1712_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1712_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1712_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1737_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1737_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1737_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1737_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1737_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1737_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2185_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2185_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2185_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2185_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2185_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2185_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2268_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2268_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2268_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2268_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2268_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2268_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2293_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2293_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2293_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2293_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2293_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2293_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2755_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2755_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2755_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2755_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2755_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2755_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2838_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2838_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2838_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2838_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2838_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2838_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2863_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2863_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2863_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2863_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2863_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2863_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3317_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3317_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3317_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3317_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3317_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3317_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3400_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3400_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3400_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3400_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3400_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3400_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3425_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3425_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3425_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3425_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3425_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3425_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3899_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3899_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3899_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3899_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3899_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3899_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3982_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3982_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3982_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3982_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3982_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3982_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4007_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4007_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4007_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4007_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4007_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4007_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4461_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4461_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4461_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4461_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4461_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4461_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4544_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4544_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4544_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4544_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4544_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4544_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4569_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4569_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4569_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4569_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4569_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4569_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_5025_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_5025_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_5025_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_5025_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_5025_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_5025_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_5108_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_5108_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_5108_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_5108_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_5108_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_5108_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_5133_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_5133_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_5133_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_5133_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_5133_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_5133_root_address : std_logic_vector(13 downto 0);
    signal arrayidx1003_3427 : std_logic_vector(31 downto 0);
    signal arrayidx1178_3901 : std_logic_vector(31 downto 0);
    signal arrayidx1221_3984 : std_logic_vector(31 downto 0);
    signal arrayidx1226_4009 : std_logic_vector(31 downto 0);
    signal arrayidx131_1157 : std_logic_vector(31 downto 0);
    signal arrayidx136_1182 : std_logic_vector(31 downto 0);
    signal arrayidx1396_4463 : std_logic_vector(31 downto 0);
    signal arrayidx1439_4546 : std_logic_vector(31 downto 0);
    signal arrayidx1444_4571 : std_logic_vector(31 downto 0);
    signal arrayidx1616_5027 : std_logic_vector(31 downto 0);
    signal arrayidx1659_5110 : std_logic_vector(31 downto 0);
    signal arrayidx1664_5135 : std_logic_vector(31 downto 0);
    signal arrayidx299_1631 : std_logic_vector(31 downto 0);
    signal arrayidx342_1714 : std_logic_vector(31 downto 0);
    signal arrayidx347_1739 : std_logic_vector(31 downto 0);
    signal arrayidx516_2187 : std_logic_vector(31 downto 0);
    signal arrayidx559_2270 : std_logic_vector(31 downto 0);
    signal arrayidx564_2295 : std_logic_vector(31 downto 0);
    signal arrayidx737_2757 : std_logic_vector(31 downto 0);
    signal arrayidx780_2840 : std_logic_vector(31 downto 0);
    signal arrayidx785_2865 : std_logic_vector(31 downto 0);
    signal arrayidx955_3319 : std_logic_vector(31 downto 0);
    signal arrayidx998_3402 : std_logic_vector(31 downto 0);
    signal arrayidx_1074 : std_logic_vector(31 downto 0);
    signal call_716 : std_logic_vector(15 downto 0);
    signal cmp1012_3451 : std_logic_vector(0 downto 0);
    signal cmp1031_3500 : std_logic_vector(0 downto 0);
    signal cmp1048_3550 : std_logic_vector(0 downto 0);
    signal cmp1127_3760 : std_logic_vector(0 downto 0);
    signal cmp1139_3798 : std_logic_vector(0 downto 0);
    signal cmp1146_3817 : std_logic_vector(0 downto 0);
    signal cmp1156_3843 : std_logic_vector(0 downto 0);
    signal cmp1235_4033 : std_logic_vector(0 downto 0);
    signal cmp1253_4076 : std_logic_vector(0 downto 0);
    signal cmp1270_4125 : std_logic_vector(0 downto 0);
    signal cmp1346_4328 : std_logic_vector(0 downto 0);
    signal cmp1356_4354 : std_logic_vector(0 downto 0);
    signal cmp1363_4373 : std_logic_vector(0 downto 0);
    signal cmp1374_4405 : std_logic_vector(0 downto 0);
    signal cmp143_1206 : std_logic_vector(0 downto 0);
    signal cmp1453_4595 : std_logic_vector(0 downto 0);
    signal cmp1472_4644 : std_logic_vector(0 downto 0);
    signal cmp1487_4682 : std_logic_vector(0 downto 0);
    signal cmp1567_4898 : std_logic_vector(0 downto 0);
    signal cmp1577_4924 : std_logic_vector(0 downto 0);
    signal cmp1584_4943 : std_logic_vector(0 downto 0);
    signal cmp1594_4969 : std_logic_vector(0 downto 0);
    signal cmp160_1255 : std_logic_vector(0 downto 0);
    signal cmp1673_5159 : std_logic_vector(0 downto 0);
    signal cmp1691_5202 : std_logic_vector(0 downto 0);
    signal cmp1706_5239 : std_logic_vector(0 downto 0);
    signal cmp176_1299 : std_logic_vector(0 downto 0);
    signal cmp249_1496 : std_logic_vector(0 downto 0);
    signal cmp260_1528 : std_logic_vector(0 downto 0);
    signal cmp267_1547 : std_logic_vector(0 downto 0);
    signal cmp277_1573 : std_logic_vector(0 downto 0);
    signal cmp356_1763 : std_logic_vector(0 downto 0);
    signal cmp374_1806 : std_logic_vector(0 downto 0);
    signal cmp390_1849 : std_logic_vector(0 downto 0);
    signal cmp465_2046 : std_logic_vector(0 downto 0);
    signal cmp476_2078 : std_logic_vector(0 downto 0);
    signal cmp483_2097 : std_logic_vector(0 downto 0);
    signal cmp494_2129 : std_logic_vector(0 downto 0);
    signal cmp56_964 : std_logic_vector(0 downto 0);
    signal cmp573_2319 : std_logic_vector(0 downto 0);
    signal cmp592_2368 : std_logic_vector(0 downto 0);
    signal cmp608_2412 : std_logic_vector(0 downto 0);
    signal cmp63_983 : std_logic_vector(0 downto 0);
    signal cmp687_2622 : std_logic_vector(0 downto 0);
    signal cmp698_2654 : std_logic_vector(0 downto 0);
    signal cmp705_2673 : std_logic_vector(0 downto 0);
    signal cmp715_2699 : std_logic_vector(0 downto 0);
    signal cmp74_1015 : std_logic_vector(0 downto 0);
    signal cmp794_2889 : std_logic_vector(0 downto 0);
    signal cmp812_2932 : std_logic_vector(0 downto 0);
    signal cmp828_2975 : std_logic_vector(0 downto 0);
    signal cmp903_3172 : std_logic_vector(0 downto 0);
    signal cmp915_3210 : std_logic_vector(0 downto 0);
    signal cmp922_3229 : std_logic_vector(0 downto 0);
    signal cmp933_3261 : std_logic_vector(0 downto 0);
    signal cmp_932 : std_logic_vector(0 downto 0);
    signal conv1008_3438 : std_logic_vector(31 downto 0);
    signal conv1023_3477 : std_logic_vector(31 downto 0);
    signal conv1025_3484 : std_logic_vector(31 downto 0);
    signal conv1025x_xlcssa_3584 : std_logic_vector(31 downto 0);
    signal conv1039_3521 : std_logic_vector(31 downto 0);
    signal conv1041_3528 : std_logic_vector(31 downto 0);
    signal conv104_896 : std_logic_vector(31 downto 0);
    signal conv1064_3596 : std_logic_vector(15 downto 0);
    signal conv1070_3606 : std_logic_vector(15 downto 0);
    signal conv1104_3646 : std_logic_vector(31 downto 0);
    signal conv1112_3661 : std_logic_vector(31 downto 0);
    signal conv1114_3676 : std_logic_vector(31 downto 0);
    signal conv1124_3753 : std_logic_vector(31 downto 0);
    signal conv1126_3685 : std_logic_vector(31 downto 0);
    signal conv1133_3774 : std_logic_vector(31 downto 0);
    signal conv1143_3810 : std_logic_vector(31 downto 0);
    signal conv1152_3831 : std_logic_vector(31 downto 0);
    signal conv1162_3855 : std_logic_vector(31 downto 0);
    signal conv1166_3860 : std_logic_vector(31 downto 0);
    signal conv1170_3700 : std_logic_vector(31 downto 0);
    signal conv1183_3913 : std_logic_vector(31 downto 0);
    signal conv1194_3726 : std_logic_vector(31 downto 0);
    signal conv1231_4020 : std_logic_vector(31 downto 0);
    signal conv1246_4059 : std_logic_vector(31 downto 0);
    signal conv1248_4066 : std_logic_vector(31 downto 0);
    signal conv1248x_xlcssa_4159 : std_logic_vector(31 downto 0);
    signal conv1261_4096 : std_logic_vector(31 downto 0);
    signal conv1263_4103 : std_logic_vector(31 downto 0);
    signal conv1288_4167 : std_logic_vector(15 downto 0);
    signal conv1323_4213 : std_logic_vector(31 downto 0);
    signal conv1331_4228 : std_logic_vector(31 downto 0);
    signal conv1333_4243 : std_logic_vector(31 downto 0);
    signal conv1343_4321 : std_logic_vector(31 downto 0);
    signal conv1345_4252 : std_logic_vector(31 downto 0);
    signal conv1352_4342 : std_logic_vector(31 downto 0);
    signal conv1360_4366 : std_logic_vector(31 downto 0);
    signal conv1369_4387 : std_logic_vector(31 downto 0);
    signal conv1380_4417 : std_logic_vector(31 downto 0);
    signal conv1384_4422 : std_logic_vector(31 downto 0);
    signal conv1388_4267 : std_logic_vector(31 downto 0);
    signal conv139_1193 : std_logic_vector(31 downto 0);
    signal conv1401_4475 : std_logic_vector(31 downto 0);
    signal conv1412_4293 : std_logic_vector(31 downto 0);
    signal conv1449_4582 : std_logic_vector(31 downto 0);
    signal conv1464_4621 : std_logic_vector(31 downto 0);
    signal conv1466_4628 : std_logic_vector(31 downto 0);
    signal conv1466x_xlcssa_4716 : std_logic_vector(31 downto 0);
    signal conv1480_4665 : std_logic_vector(31 downto 0);
    signal conv1482_4672 : std_logic_vector(31 downto 0);
    signal conv1503_4728 : std_logic_vector(15 downto 0);
    signal conv1509_4738 : std_logic_vector(15 downto 0);
    signal conv153_1232 : std_logic_vector(31 downto 0);
    signal conv1544_4784 : std_logic_vector(31 downto 0);
    signal conv1552_4799 : std_logic_vector(31 downto 0);
    signal conv1554_4814 : std_logic_vector(31 downto 0);
    signal conv155_1239 : std_logic_vector(31 downto 0);
    signal conv155x_xlcssa_1329 : std_logic_vector(31 downto 0);
    signal conv1564_4891 : std_logic_vector(31 downto 0);
    signal conv1566_4823 : std_logic_vector(31 downto 0);
    signal conv1573_4912 : std_logic_vector(31 downto 0);
    signal conv1581_4936 : std_logic_vector(31 downto 0);
    signal conv1590_4957 : std_logic_vector(31 downto 0);
    signal conv1600_4981 : std_logic_vector(31 downto 0);
    signal conv1604_4986 : std_logic_vector(31 downto 0);
    signal conv1608_4838 : std_logic_vector(31 downto 0);
    signal conv1621_5039 : std_logic_vector(31 downto 0);
    signal conv1632_4864 : std_logic_vector(31 downto 0);
    signal conv1669_5146 : std_logic_vector(31 downto 0);
    signal conv1684_5185 : std_logic_vector(31 downto 0);
    signal conv1686_5192 : std_logic_vector(31 downto 0);
    signal conv168_1276 : std_logic_vector(31 downto 0);
    signal conv1699_5222 : std_logic_vector(31 downto 0);
    signal conv1701_5229 : std_logic_vector(31 downto 0);
    signal conv170_1283 : std_logic_vector(31 downto 0);
    signal conv190_1341 : std_logic_vector(15 downto 0);
    signal conv226_1381 : std_logic_vector(31 downto 0);
    signal conv234_1396 : std_logic_vector(31 downto 0);
    signal conv236_1411 : std_logic_vector(31 downto 0);
    signal conv246_1489 : std_logic_vector(31 downto 0);
    signal conv248_1420 : std_logic_vector(31 downto 0);
    signal conv255_1510 : std_logic_vector(31 downto 0);
    signal conv264_1540 : std_logic_vector(31 downto 0);
    signal conv273_1561 : std_logic_vector(31 downto 0);
    signal conv283_1585 : std_logic_vector(31 downto 0);
    signal conv287_1590 : std_logic_vector(31 downto 0);
    signal conv291_1435 : std_logic_vector(31 downto 0);
    signal conv2_751 : std_logic_vector(7 downto 0);
    signal conv304_1643 : std_logic_vector(31 downto 0);
    signal conv315_1461 : std_logic_vector(31 downto 0);
    signal conv31_811 : std_logic_vector(31 downto 0);
    signal conv33_815 : std_logic_vector(31 downto 0);
    signal conv352_1750 : std_logic_vector(31 downto 0);
    signal conv367_1789 : std_logic_vector(31 downto 0);
    signal conv369_1796 : std_logic_vector(31 downto 0);
    signal conv369x_xlcssa_1883 : std_logic_vector(31 downto 0);
    signal conv37_831 : std_logic_vector(31 downto 0);
    signal conv382_1826 : std_logic_vector(31 downto 0);
    signal conv384_1833 : std_logic_vector(31 downto 0);
    signal conv39_846 : std_logic_vector(31 downto 0);
    signal conv408_1891 : std_logic_vector(15 downto 0);
    signal conv442_1931 : std_logic_vector(31 downto 0);
    signal conv450_1946 : std_logic_vector(31 downto 0);
    signal conv452_1961 : std_logic_vector(31 downto 0);
    signal conv462_2039 : std_logic_vector(31 downto 0);
    signal conv464_1970 : std_logic_vector(31 downto 0);
    signal conv46_925 : std_logic_vector(31 downto 0);
    signal conv471_2060 : std_logic_vector(31 downto 0);
    signal conv480_2090 : std_logic_vector(31 downto 0);
    signal conv489_2111 : std_logic_vector(31 downto 0);
    signal conv48_855 : std_logic_vector(31 downto 0);
    signal conv4_770 : std_logic_vector(7 downto 0);
    signal conv500_2141 : std_logic_vector(31 downto 0);
    signal conv504_2146 : std_logic_vector(31 downto 0);
    signal conv508_1985 : std_logic_vector(31 downto 0);
    signal conv521_2199 : std_logic_vector(31 downto 0);
    signal conv532_2011 : std_logic_vector(31 downto 0);
    signal conv53_946 : std_logic_vector(31 downto 0);
    signal conv569_2306 : std_logic_vector(31 downto 0);
    signal conv584_2345 : std_logic_vector(31 downto 0);
    signal conv586_2352 : std_logic_vector(31 downto 0);
    signal conv586x_xlcssa_2446 : std_logic_vector(31 downto 0);
    signal conv600_2389 : std_logic_vector(31 downto 0);
    signal conv602_2396 : std_logic_vector(31 downto 0);
    signal conv60_976 : std_logic_vector(31 downto 0);
    signal conv624_2458 : std_logic_vector(15 downto 0);
    signal conv630_2468 : std_logic_vector(15 downto 0);
    signal conv664_2508 : std_logic_vector(31 downto 0);
    signal conv672_2523 : std_logic_vector(31 downto 0);
    signal conv674_2538 : std_logic_vector(31 downto 0);
    signal conv684_2615 : std_logic_vector(31 downto 0);
    signal conv686_2547 : std_logic_vector(31 downto 0);
    signal conv693_2636 : std_logic_vector(31 downto 0);
    signal conv69_997 : std_logic_vector(31 downto 0);
    signal conv702_2666 : std_logic_vector(31 downto 0);
    signal conv711_2687 : std_logic_vector(31 downto 0);
    signal conv721_2711 : std_logic_vector(31 downto 0);
    signal conv725_2716 : std_logic_vector(31 downto 0);
    signal conv729_2562 : std_logic_vector(31 downto 0);
    signal conv742_2769 : std_logic_vector(31 downto 0);
    signal conv753_2588 : std_logic_vector(31 downto 0);
    signal conv78_1027 : std_logic_vector(31 downto 0);
    signal conv790_2876 : std_logic_vector(31 downto 0);
    signal conv805_2915 : std_logic_vector(31 downto 0);
    signal conv807_2922 : std_logic_vector(31 downto 0);
    signal conv807x_xlcssa_3009 : std_logic_vector(31 downto 0);
    signal conv820_2952 : std_logic_vector(31 downto 0);
    signal conv822_2959 : std_logic_vector(31 downto 0);
    signal conv82_1032 : std_logic_vector(31 downto 0);
    signal conv846_3017 : std_logic_vector(15 downto 0);
    signal conv86_870 : std_logic_vector(31 downto 0);
    signal conv880_3057 : std_logic_vector(31 downto 0);
    signal conv888_3072 : std_logic_vector(31 downto 0);
    signal conv890_3087 : std_logic_vector(31 downto 0);
    signal conv900_3165 : std_logic_vector(31 downto 0);
    signal conv902_3096 : std_logic_vector(31 downto 0);
    signal conv909_3186 : std_logic_vector(31 downto 0);
    signal conv919_3222 : std_logic_vector(31 downto 0);
    signal conv928_3243 : std_logic_vector(31 downto 0);
    signal conv939_3273 : std_logic_vector(31 downto 0);
    signal conv943_3278 : std_logic_vector(31 downto 0);
    signal conv947_3111 : std_logic_vector(31 downto 0);
    signal conv94_1086 : std_logic_vector(31 downto 0);
    signal conv960_3331 : std_logic_vector(31 downto 0);
    signal conv971_3137 : std_logic_vector(31 downto 0);
    signal conv_732 : std_logic_vector(7 downto 0);
    signal div1026_3490 : std_logic_vector(31 downto 0);
    signal div1043_3540 : std_logic_vector(31 downto 0);
    signal div1065_3602 : std_logic_vector(15 downto 0);
    signal div1071_3612 : std_logic_vector(15 downto 0);
    signal div1135_3786 : std_logic_vector(31 downto 0);
    signal div1265_4115 : std_logic_vector(31 downto 0);
    signal div1289_4173 : std_logic_vector(15 downto 0);
    signal div1370_4393 : std_logic_vector(31 downto 0);
    signal div1467_4634 : std_logic_vector(31 downto 0);
    signal div1504_4734 : std_logic_vector(15 downto 0);
    signal div1511_4750 : std_logic_vector(15 downto 0);
    signal div156_1245 : std_logic_vector(31 downto 0);
    signal div171_1289 : std_logic_vector(31 downto 0);
    signal div191_1347 : std_logic_vector(15 downto 0);
    signal div256_1516 : std_logic_vector(31 downto 0);
    signal div385_1839 : std_logic_vector(31 downto 0);
    signal div409_1897 : std_logic_vector(15 downto 0);
    signal div472_2066 : std_logic_vector(31 downto 0);
    signal div490_2117 : std_logic_vector(31 downto 0);
    signal div587_2358 : std_logic_vector(31 downto 0);
    signal div603_2402 : std_logic_vector(31 downto 0);
    signal div625_2464 : std_logic_vector(15 downto 0);
    signal div631_2474 : std_logic_vector(15 downto 0);
    signal div694_2642 : std_logic_vector(31 downto 0);
    signal div70_1003 : std_logic_vector(31 downto 0);
    signal div823_2965 : std_logic_vector(31 downto 0);
    signal div847_3023 : std_logic_vector(15 downto 0);
    signal div911_3198 : std_logic_vector(31 downto 0);
    signal div929_3249 : std_logic_vector(31 downto 0);
    signal div_952 : std_logic_vector(31 downto 0);
    signal i1068x_x1x_xph_4140 : std_logic_vector(15 downto 0);
    signal i1068x_x2_3736 : std_logic_vector(15 downto 0);
    signal i1286x_x1x_xph_4697 : std_logic_vector(15 downto 0);
    signal i1286x_x2_4303 : std_logic_vector(15 downto 0);
    signal i1507x_x1x_xph_5254 : std_logic_vector(15 downto 0);
    signal i1507x_x2_4874 : std_logic_vector(15 downto 0);
    signal i194x_x1x_xph_1863 : std_logic_vector(15 downto 0);
    signal i194x_x2_1470 : std_logic_vector(15 downto 0);
    signal i406x_x1x_xph_2427 : std_logic_vector(15 downto 0);
    signal i406x_x2_2021 : std_logic_vector(15 downto 0);
    signal i628x_x1x_xph_2990 : std_logic_vector(15 downto 0);
    signal i628x_x2_2598 : std_logic_vector(15 downto 0);
    signal i844x_x1x_xph_3565 : std_logic_vector(15 downto 0);
    signal i844x_x2_3147 : std_logic_vector(15 downto 0);
    signal iNsTr_0_724 : std_logic_vector(31 downto 0);
    signal iNsTr_101_4193 : std_logic_vector(31 downto 0);
    signal iNsTr_102_4205 : std_logic_vector(31 downto 0);
    signal iNsTr_117_4764 : std_logic_vector(31 downto 0);
    signal iNsTr_118_4776 : std_logic_vector(31 downto 0);
    signal iNsTr_21_1361 : std_logic_vector(31 downto 0);
    signal iNsTr_22_1373 : std_logic_vector(31 downto 0);
    signal iNsTr_2_743 : std_logic_vector(31 downto 0);
    signal iNsTr_37_1911 : std_logic_vector(31 downto 0);
    signal iNsTr_38_1923 : std_logic_vector(31 downto 0);
    signal iNsTr_4_762 : std_logic_vector(31 downto 0);
    signal iNsTr_53_2488 : std_logic_vector(31 downto 0);
    signal iNsTr_54_2500 : std_logic_vector(31 downto 0);
    signal iNsTr_69_3037 : std_logic_vector(31 downto 0);
    signal iNsTr_70_3049 : std_logic_vector(31 downto 0);
    signal iNsTr_7_791 : std_logic_vector(31 downto 0);
    signal iNsTr_85_3626 : std_logic_vector(31 downto 0);
    signal iNsTr_86_3638 : std_logic_vector(31 downto 0);
    signal iNsTr_8_803 : std_logic_vector(31 downto 0);
    signal idxprom1002_3420 : std_logic_vector(63 downto 0);
    signal idxprom1177_3894 : std_logic_vector(63 downto 0);
    signal idxprom1220_3977 : std_logic_vector(63 downto 0);
    signal idxprom1225_4002 : std_logic_vector(63 downto 0);
    signal idxprom130_1150 : std_logic_vector(63 downto 0);
    signal idxprom135_1175 : std_logic_vector(63 downto 0);
    signal idxprom1395_4456 : std_logic_vector(63 downto 0);
    signal idxprom1438_4539 : std_logic_vector(63 downto 0);
    signal idxprom1443_4564 : std_logic_vector(63 downto 0);
    signal idxprom1615_5020 : std_logic_vector(63 downto 0);
    signal idxprom1658_5103 : std_logic_vector(63 downto 0);
    signal idxprom1663_5128 : std_logic_vector(63 downto 0);
    signal idxprom298_1624 : std_logic_vector(63 downto 0);
    signal idxprom341_1707 : std_logic_vector(63 downto 0);
    signal idxprom346_1732 : std_logic_vector(63 downto 0);
    signal idxprom515_2180 : std_logic_vector(63 downto 0);
    signal idxprom558_2263 : std_logic_vector(63 downto 0);
    signal idxprom563_2288 : std_logic_vector(63 downto 0);
    signal idxprom736_2750 : std_logic_vector(63 downto 0);
    signal idxprom779_2833 : std_logic_vector(63 downto 0);
    signal idxprom784_2858 : std_logic_vector(63 downto 0);
    signal idxprom954_3312 : std_logic_vector(63 downto 0);
    signal idxprom997_3395 : std_logic_vector(63 downto 0);
    signal idxprom_1067 : std_logic_vector(63 downto 0);
    signal inc1021_3472 : std_logic_vector(15 downto 0);
    signal inc1036_3504 : std_logic_vector(15 downto 0);
    signal inc1036x_xi844x_x2_3509 : std_logic_vector(15 downto 0);
    signal inc1244_4054 : std_logic_vector(15 downto 0);
    signal inc1258_4080 : std_logic_vector(15 downto 0);
    signal inc1258x_xi1068x_x2_4085 : std_logic_vector(15 downto 0);
    signal inc1462_4616 : std_logic_vector(15 downto 0);
    signal inc1477_4648 : std_logic_vector(15 downto 0);
    signal inc1477x_xi1286x_x2_4653 : std_logic_vector(15 downto 0);
    signal inc165_1259 : std_logic_vector(15 downto 0);
    signal inc165x_xix_x2_1264 : std_logic_vector(15 downto 0);
    signal inc1682_5180 : std_logic_vector(15 downto 0);
    signal inc1696_5206 : std_logic_vector(15 downto 0);
    signal inc1696x_xi1507x_x2_5211 : std_logic_vector(15 downto 0);
    signal inc365_1784 : std_logic_vector(15 downto 0);
    signal inc379_1810 : std_logic_vector(15 downto 0);
    signal inc379x_xi194x_x2_1815 : std_logic_vector(15 downto 0);
    signal inc582_2340 : std_logic_vector(15 downto 0);
    signal inc597_2372 : std_logic_vector(15 downto 0);
    signal inc597x_xi406x_x2_2377 : std_logic_vector(15 downto 0);
    signal inc803_2910 : std_logic_vector(15 downto 0);
    signal inc817_2936 : std_logic_vector(15 downto 0);
    signal inc817x_xi628x_x2_2941 : std_logic_vector(15 downto 0);
    signal inc_1227 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_1313 : std_logic_vector(15 downto 0);
    signal ix_x2_906 : std_logic_vector(15 downto 0);
    signal j1118x_x0x_xph_4146 : std_logic_vector(15 downto 0);
    signal j1118x_x1_3742 : std_logic_vector(15 downto 0);
    signal j1118x_x2_4091 : std_logic_vector(15 downto 0);
    signal j1337x_x0x_xph_4703 : std_logic_vector(15 downto 0);
    signal j1337x_x1_4309 : std_logic_vector(15 downto 0);
    signal j1337x_x2_4660 : std_logic_vector(15 downto 0);
    signal j1558x_x0x_xph_5260 : std_logic_vector(15 downto 0);
    signal j1558x_x1_4880 : std_logic_vector(15 downto 0);
    signal j1558x_x2_5217 : std_logic_vector(15 downto 0);
    signal j240x_x0x_xph_1857 : std_logic_vector(15 downto 0);
    signal j240x_x1_1464 : std_logic_vector(15 downto 0);
    signal j240x_x2_1821 : std_logic_vector(15 downto 0);
    signal j456x_x0x_xph_2433 : std_logic_vector(15 downto 0);
    signal j456x_x1_2027 : std_logic_vector(15 downto 0);
    signal j456x_x2_2384 : std_logic_vector(15 downto 0);
    signal j678x_x0x_xph_2996 : std_logic_vector(15 downto 0);
    signal j678x_x1_2604 : std_logic_vector(15 downto 0);
    signal j678x_x2_2947 : std_logic_vector(15 downto 0);
    signal j894x_x0x_xph_3571 : std_logic_vector(15 downto 0);
    signal j894x_x1_3153 : std_logic_vector(15 downto 0);
    signal j894x_x2_3516 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_1307 : std_logic_vector(15 downto 0);
    signal jx_x1_899 : std_logic_vector(15 downto 0);
    signal jx_x2_1271 : std_logic_vector(15 downto 0);
    signal k1060x_x0x_xph_4133 : std_logic_vector(15 downto 0);
    signal k1060x_x1_3729 : std_logic_vector(15 downto 0);
    signal k1282x_x0x_xph_4690 : std_logic_vector(15 downto 0);
    signal k1282x_x1_4296 : std_logic_vector(15 downto 0);
    signal k1499x_x0x_xph_5247 : std_logic_vector(15 downto 0);
    signal k1499x_x1_4867 : std_logic_vector(15 downto 0);
    signal k186x_x0x_xph_1869 : std_logic_vector(15 downto 0);
    signal k186x_x1_1477 : std_logic_vector(15 downto 0);
    signal k402x_x0x_xph_2420 : std_logic_vector(15 downto 0);
    signal k402x_x1_2014 : std_logic_vector(15 downto 0);
    signal k620x_x0x_xph_2983 : std_logic_vector(15 downto 0);
    signal k620x_x1_2591 : std_logic_vector(15 downto 0);
    signal k840x_x0x_xph_3558 : std_logic_vector(15 downto 0);
    signal k840x_x1_3140 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_1319 : std_logic_vector(15 downto 0);
    signal kx_x1_913 : std_logic_vector(15 downto 0);
    signal mul101_1096 : std_logic_vector(31 downto 0);
    signal mul1042_3534 : std_logic_vector(31 downto 0);
    signal mul1107_3712 : std_logic_vector(31 downto 0);
    signal mul110_1106 : std_logic_vector(31 downto 0);
    signal mul1115_3681 : std_logic_vector(31 downto 0);
    signal mul1134_3780 : std_logic_vector(31 downto 0);
    signal mul1167_3865 : std_logic_vector(31 downto 0);
    signal mul1173_3870 : std_logic_vector(31 downto 0);
    signal mul1191_3923 : std_logic_vector(31 downto 0);
    signal mul1200_3933 : std_logic_vector(31 downto 0);
    signal mul120_1121 : std_logic_vector(31 downto 0);
    signal mul1210_3948 : std_logic_vector(31 downto 0);
    signal mul1216_3953 : std_logic_vector(31 downto 0);
    signal mul1264_4109 : std_logic_vector(31 downto 0);
    signal mul126_1126 : std_logic_vector(31 downto 0);
    signal mul1290_4179 : std_logic_vector(15 downto 0);
    signal mul1326_4279 : std_logic_vector(31 downto 0);
    signal mul1334_4248 : std_logic_vector(31 downto 0);
    signal mul1385_4427 : std_logic_vector(31 downto 0);
    signal mul1391_4432 : std_logic_vector(31 downto 0);
    signal mul1409_4485 : std_logic_vector(31 downto 0);
    signal mul1418_4495 : std_logic_vector(31 downto 0);
    signal mul1428_4510 : std_logic_vector(31 downto 0);
    signal mul1434_4515 : std_logic_vector(31 downto 0);
    signal mul1510_4744 : std_logic_vector(15 downto 0);
    signal mul1547_4850 : std_logic_vector(31 downto 0);
    signal mul1555_4819 : std_logic_vector(31 downto 0);
    signal mul1605_4991 : std_logic_vector(31 downto 0);
    signal mul1611_4996 : std_logic_vector(31 downto 0);
    signal mul1629_5049 : std_logic_vector(31 downto 0);
    signal mul1638_5059 : std_logic_vector(31 downto 0);
    signal mul1648_5074 : std_logic_vector(31 downto 0);
    signal mul1654_5079 : std_logic_vector(31 downto 0);
    signal mul229_1447 : std_logic_vector(31 downto 0);
    signal mul237_1416 : std_logic_vector(31 downto 0);
    signal mul288_1595 : std_logic_vector(31 downto 0);
    signal mul294_1600 : std_logic_vector(31 downto 0);
    signal mul312_1653 : std_logic_vector(31 downto 0);
    signal mul321_1663 : std_logic_vector(31 downto 0);
    signal mul331_1678 : std_logic_vector(31 downto 0);
    signal mul337_1683 : std_logic_vector(31 downto 0);
    signal mul40_851 : std_logic_vector(31 downto 0);
    signal mul445_1997 : std_logic_vector(31 downto 0);
    signal mul453_1966 : std_logic_vector(31 downto 0);
    signal mul505_2151 : std_logic_vector(31 downto 0);
    signal mul511_2156 : std_logic_vector(31 downto 0);
    signal mul529_2209 : std_logic_vector(31 downto 0);
    signal mul538_2219 : std_logic_vector(31 downto 0);
    signal mul548_2234 : std_logic_vector(31 downto 0);
    signal mul554_2239 : std_logic_vector(31 downto 0);
    signal mul667_2574 : std_logic_vector(31 downto 0);
    signal mul675_2543 : std_logic_vector(31 downto 0);
    signal mul726_2721 : std_logic_vector(31 downto 0);
    signal mul732_2726 : std_logic_vector(31 downto 0);
    signal mul750_2779 : std_logic_vector(31 downto 0);
    signal mul759_2789 : std_logic_vector(31 downto 0);
    signal mul769_2804 : std_logic_vector(31 downto 0);
    signal mul775_2809 : std_logic_vector(31 downto 0);
    signal mul83_1037 : std_logic_vector(31 downto 0);
    signal mul883_3123 : std_logic_vector(31 downto 0);
    signal mul891_3092 : std_logic_vector(31 downto 0);
    signal mul89_1042 : std_logic_vector(31 downto 0);
    signal mul910_3192 : std_logic_vector(31 downto 0);
    signal mul944_3283 : std_logic_vector(31 downto 0);
    signal mul950_3288 : std_logic_vector(31 downto 0);
    signal mul968_3341 : std_logic_vector(31 downto 0);
    signal mul977_3351 : std_logic_vector(31 downto 0);
    signal mul987_3366 : std_logic_vector(31 downto 0);
    signal mul993_3371 : std_logic_vector(31 downto 0);
    signal mul_882 : std_logic_vector(31 downto 0);
    signal ptr_deref_1076_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1076_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1076_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1076_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1076_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1076_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1160_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1160_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1160_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1160_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1160_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1184_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1184_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1184_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1184_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1184_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1184_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1364_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1364_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1364_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1364_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1364_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1376_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1376_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1376_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1376_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1376_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1633_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1633_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1633_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1633_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1633_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1633_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1717_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1717_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1717_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1717_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1717_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1741_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1741_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1741_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1741_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1741_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1741_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1914_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1914_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1914_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1914_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1914_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1926_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1926_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1926_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1926_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1926_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2189_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2189_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2189_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2189_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2189_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2189_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2273_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2273_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2273_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2273_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2273_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2297_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2297_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2297_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2297_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2297_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2297_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2491_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2491_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2491_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2491_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2491_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2503_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2503_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2503_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2503_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2503_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2759_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2759_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2759_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2759_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2759_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2759_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2843_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2843_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2843_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2843_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2843_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2867_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2867_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2867_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2867_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2867_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2867_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3040_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3040_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3040_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3040_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3040_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3052_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3052_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3052_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3052_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3052_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3321_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3321_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3321_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3321_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3321_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3321_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3405_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3405_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3405_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3405_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3405_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3429_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3429_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3429_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3429_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3429_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3429_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3629_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3629_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3629_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3629_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3629_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3641_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3641_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3641_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3641_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3641_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3903_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3903_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3903_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3903_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3903_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3903_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3987_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3987_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3987_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3987_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3987_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4011_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4011_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4011_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4011_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4011_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4011_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4196_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_4196_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4196_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4196_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4196_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4208_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_4208_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4208_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4208_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4208_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4465_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4465_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4465_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4465_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4465_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4465_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4549_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4549_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4549_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4549_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4549_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4573_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4573_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4573_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4573_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4573_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4573_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4767_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_4767_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4767_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4767_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4767_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4779_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_4779_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4779_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4779_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4779_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_5029_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_5029_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_5029_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_5029_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_5029_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_5029_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_5113_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_5113_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_5113_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_5113_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_5113_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_5137_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_5137_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_5137_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_5137_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_5137_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_5137_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_727_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_727_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_727_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_727_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_727_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_746_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_746_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_746_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_746_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_746_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_765_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_765_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_765_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_765_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_765_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_794_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_794_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_794_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_794_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_794_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_806_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_806_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_806_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_806_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_806_word_offset_0 : std_logic_vector(6 downto 0);
    signal sext1717_887 : std_logic_vector(31 downto 0);
    signal sext1718_1402 : std_logic_vector(31 downto 0);
    signal sext1719_1452 : std_logic_vector(31 downto 0);
    signal sext1720_1952 : std_logic_vector(31 downto 0);
    signal sext1721_2002 : std_logic_vector(31 downto 0);
    signal sext1722_2529 : std_logic_vector(31 downto 0);
    signal sext1723_2579 : std_logic_vector(31 downto 0);
    signal sext1724_3078 : std_logic_vector(31 downto 0);
    signal sext1725_3128 : std_logic_vector(31 downto 0);
    signal sext1726_3667 : std_logic_vector(31 downto 0);
    signal sext1727_3717 : std_logic_vector(31 downto 0);
    signal sext1728_4234 : std_logic_vector(31 downto 0);
    signal sext1729_4284 : std_logic_vector(31 downto 0);
    signal sext1730_4805 : std_logic_vector(31 downto 0);
    signal sext1731_4855 : std_logic_vector(31 downto 0);
    signal sext1764_821 : std_logic_vector(31 downto 0);
    signal sext1765_861 : std_logic_vector(31 downto 0);
    signal sext1766_1387 : std_logic_vector(31 downto 0);
    signal sext1767_1426 : std_logic_vector(31 downto 0);
    signal sext1768_1937 : std_logic_vector(31 downto 0);
    signal sext1769_1976 : std_logic_vector(31 downto 0);
    signal sext1770_2514 : std_logic_vector(31 downto 0);
    signal sext1771_2553 : std_logic_vector(31 downto 0);
    signal sext1772_3063 : std_logic_vector(31 downto 0);
    signal sext1773_3102 : std_logic_vector(31 downto 0);
    signal sext1774_3652 : std_logic_vector(31 downto 0);
    signal sext1775_3691 : std_logic_vector(31 downto 0);
    signal sext1776_4219 : std_logic_vector(31 downto 0);
    signal sext1777_4258 : std_logic_vector(31 downto 0);
    signal sext1778_4790 : std_logic_vector(31 downto 0);
    signal sext1779_4829 : std_logic_vector(31 downto 0);
    signal sext_837 : std_logic_vector(31 downto 0);
    signal shl1029_3117 : std_logic_vector(31 downto 0);
    signal shl1251_3706 : std_logic_vector(31 downto 0);
    signal shl1470_4273 : std_logic_vector(31 downto 0);
    signal shl1689_4844 : std_logic_vector(31 downto 0);
    signal shl372_1441 : std_logic_vector(31 downto 0);
    signal shl590_1991 : std_logic_vector(31 downto 0);
    signal shl810_2568 : std_logic_vector(31 downto 0);
    signal shl_876 : std_logic_vector(31 downto 0);
    signal shr1001_3415 : std_logic_vector(31 downto 0);
    signal shr1176_3889 : std_logic_vector(31 downto 0);
    signal shr1219_3972 : std_logic_vector(31 downto 0);
    signal shr1224_3997 : std_logic_vector(31 downto 0);
    signal shr129_1145 : std_logic_vector(31 downto 0);
    signal shr134_1170 : std_logic_vector(31 downto 0);
    signal shr1394_4451 : std_logic_vector(31 downto 0);
    signal shr1437_4534 : std_logic_vector(31 downto 0);
    signal shr1442_4559 : std_logic_vector(31 downto 0);
    signal shr1614_5015 : std_logic_vector(31 downto 0);
    signal shr1657_5098 : std_logic_vector(31 downto 0);
    signal shr1662_5123 : std_logic_vector(31 downto 0);
    signal shr297_1619 : std_logic_vector(31 downto 0);
    signal shr340_1702 : std_logic_vector(31 downto 0);
    signal shr345_1727 : std_logic_vector(31 downto 0);
    signal shr514_2175 : std_logic_vector(31 downto 0);
    signal shr557_2258 : std_logic_vector(31 downto 0);
    signal shr562_2283 : std_logic_vector(31 downto 0);
    signal shr735_2745 : std_logic_vector(31 downto 0);
    signal shr778_2828 : std_logic_vector(31 downto 0);
    signal shr783_2853 : std_logic_vector(31 downto 0);
    signal shr953_3307 : std_logic_vector(31 downto 0);
    signal shr996_3390 : std_logic_vector(31 downto 0);
    signal shr_1061 : std_logic_vector(31 downto 0);
    signal sub109_1101 : std_logic_vector(31 downto 0);
    signal sub1190_3918 : std_logic_vector(31 downto 0);
    signal sub1199_3928 : std_logic_vector(31 downto 0);
    signal sub1408_4480 : std_logic_vector(31 downto 0);
    signal sub1417_4490 : std_logic_vector(31 downto 0);
    signal sub1628_5044 : std_logic_vector(31 downto 0);
    signal sub1637_5054 : std_logic_vector(31 downto 0);
    signal sub311_1648 : std_logic_vector(31 downto 0);
    signal sub320_1658 : std_logic_vector(31 downto 0);
    signal sub528_2204 : std_logic_vector(31 downto 0);
    signal sub537_2214 : std_logic_vector(31 downto 0);
    signal sub749_2774 : std_logic_vector(31 downto 0);
    signal sub758_2784 : std_logic_vector(31 downto 0);
    signal sub967_3336 : std_logic_vector(31 downto 0);
    signal sub976_3346 : std_logic_vector(31 downto 0);
    signal sub_1091 : std_logic_vector(31 downto 0);
    signal tmp1024_3480 : std_logic_vector(7 downto 0);
    signal tmp1024x_xlcssa_3588 : std_logic_vector(7 downto 0);
    signal tmp1040_3524 : std_logic_vector(7 downto 0);
    signal tmp1040x_xlcssa_3580 : std_logic_vector(7 downto 0);
    signal tmp1075_3615 : std_logic_vector(7 downto 0);
    signal tmp1079_3618 : std_logic_vector(7 downto 0);
    signal tmp1091_3630 : std_logic_vector(31 downto 0);
    signal tmp1095_3642 : std_logic_vector(31 downto 0);
    signal tmp1132_3770 : std_logic_vector(7 downto 0);
    signal tmp1151_3827 : std_logic_vector(7 downto 0);
    signal tmp1222_3988 : std_logic_vector(63 downto 0);
    signal tmp1247_4062 : std_logic_vector(7 downto 0);
    signal tmp1262_4099 : std_logic_vector(7 downto 0);
    signal tmp1262x_xlcssa_4155 : std_logic_vector(7 downto 0);
    signal tmp1294_4182 : std_logic_vector(7 downto 0);
    signal tmp1298_4185 : std_logic_vector(7 downto 0);
    signal tmp12_780 : std_logic_vector(7 downto 0);
    signal tmp1310_4197 : std_logic_vector(31 downto 0);
    signal tmp1314_4209 : std_logic_vector(31 downto 0);
    signal tmp132_1161 : std_logic_vector(63 downto 0);
    signal tmp1351_4338 : std_logic_vector(7 downto 0);
    signal tmp1368_4383 : std_logic_vector(7 downto 0);
    signal tmp1440_4550 : std_logic_vector(63 downto 0);
    signal tmp1465_4624 : std_logic_vector(7 downto 0);
    signal tmp1465x_xlcssa_4720 : std_logic_vector(7 downto 0);
    signal tmp1481_4668 : std_logic_vector(7 downto 0);
    signal tmp1481x_xlcssa_4712 : std_logic_vector(7 downto 0);
    signal tmp1515_4753 : std_logic_vector(7 downto 0);
    signal tmp1519_4756 : std_logic_vector(7 downto 0);
    signal tmp1531_4768 : std_logic_vector(31 downto 0);
    signal tmp1535_4780 : std_logic_vector(31 downto 0);
    signal tmp154_1235 : std_logic_vector(7 downto 0);
    signal tmp154x_xlcssa_1333 : std_logic_vector(7 downto 0);
    signal tmp1572_4908 : std_logic_vector(7 downto 0);
    signal tmp1589_4953 : std_logic_vector(7 downto 0);
    signal tmp15_783 : std_logic_vector(7 downto 0);
    signal tmp1660_5114 : std_logic_vector(63 downto 0);
    signal tmp1685_5188 : std_logic_vector(7 downto 0);
    signal tmp169_1279 : std_logic_vector(7 downto 0);
    signal tmp1700_5225 : std_logic_vector(7 downto 0);
    signal tmp197_1350 : std_logic_vector(7 downto 0);
    signal tmp1_747 : std_logic_vector(31 downto 0);
    signal tmp201_1353 : std_logic_vector(7 downto 0);
    signal tmp213_1365 : std_logic_vector(31 downto 0);
    signal tmp217_1377 : std_logic_vector(31 downto 0);
    signal tmp21_795 : std_logic_vector(31 downto 0);
    signal tmp24_807 : std_logic_vector(31 downto 0);
    signal tmp254_1506 : std_logic_vector(7 downto 0);
    signal tmp272_1557 : std_logic_vector(7 downto 0);
    signal tmp343_1718 : std_logic_vector(63 downto 0);
    signal tmp368_1792 : std_logic_vector(7 downto 0);
    signal tmp383_1829 : std_logic_vector(7 downto 0);
    signal tmp383x_xlcssa_1879 : std_logic_vector(7 downto 0);
    signal tmp3_766 : std_logic_vector(31 downto 0);
    signal tmp413_1900 : std_logic_vector(7 downto 0);
    signal tmp417_1903 : std_logic_vector(7 downto 0);
    signal tmp429_1915 : std_logic_vector(31 downto 0);
    signal tmp433_1927 : std_logic_vector(31 downto 0);
    signal tmp470_2056 : std_logic_vector(7 downto 0);
    signal tmp488_2107 : std_logic_vector(7 downto 0);
    signal tmp52_942 : std_logic_vector(7 downto 0);
    signal tmp560_2274 : std_logic_vector(63 downto 0);
    signal tmp585_2348 : std_logic_vector(7 downto 0);
    signal tmp585x_xlcssa_2450 : std_logic_vector(7 downto 0);
    signal tmp601_2392 : std_logic_vector(7 downto 0);
    signal tmp601x_xlcssa_2442 : std_logic_vector(7 downto 0);
    signal tmp635_2477 : std_logic_vector(7 downto 0);
    signal tmp639_2480 : std_logic_vector(7 downto 0);
    signal tmp651_2492 : std_logic_vector(31 downto 0);
    signal tmp655_2504 : std_logic_vector(31 downto 0);
    signal tmp68_993 : std_logic_vector(7 downto 0);
    signal tmp692_2632 : std_logic_vector(7 downto 0);
    signal tmp710_2683 : std_logic_vector(7 downto 0);
    signal tmp781_2844 : std_logic_vector(63 downto 0);
    signal tmp806_2918 : std_logic_vector(7 downto 0);
    signal tmp821_2955 : std_logic_vector(7 downto 0);
    signal tmp821x_xlcssa_3005 : std_logic_vector(7 downto 0);
    signal tmp851_3026 : std_logic_vector(7 downto 0);
    signal tmp855_3029 : std_logic_vector(7 downto 0);
    signal tmp867_3041 : std_logic_vector(31 downto 0);
    signal tmp871_3053 : std_logic_vector(31 downto 0);
    signal tmp908_3182 : std_logic_vector(7 downto 0);
    signal tmp927_3239 : std_logic_vector(7 downto 0);
    signal tmp999_3406 : std_logic_vector(63 downto 0);
    signal tmp9_777 : std_logic_vector(7 downto 0);
    signal tmp_728 : std_logic_vector(31 downto 0);
    signal type_cast_1001_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1011_wire : std_logic_vector(31 downto 0);
    signal type_cast_1013_wire : std_logic_vector(31 downto 0);
    signal type_cast_1025_wire : std_logic_vector(31 downto 0);
    signal type_cast_1030_wire : std_logic_vector(31 downto 0);
    signal type_cast_1055_wire : std_logic_vector(31 downto 0);
    signal type_cast_1058_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1065_wire : std_logic_vector(63 downto 0);
    signal type_cast_1078_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1084_wire : std_logic_vector(31 downto 0);
    signal type_cast_1139_wire : std_logic_vector(31 downto 0);
    signal type_cast_1142_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1148_wire : std_logic_vector(63 downto 0);
    signal type_cast_1164_wire : std_logic_vector(31 downto 0);
    signal type_cast_1167_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1173_wire : std_logic_vector(63 downto 0);
    signal type_cast_1191_wire : std_logic_vector(31 downto 0);
    signal type_cast_1197_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1202_wire : std_logic_vector(31 downto 0);
    signal type_cast_1204_wire : std_logic_vector(31 downto 0);
    signal type_cast_1217_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1225_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1230_wire : std_logic_vector(31 downto 0);
    signal type_cast_1243_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1268_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1274_wire : std_logic_vector(31 downto 0);
    signal type_cast_1287_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1310_wire : std_logic_vector(15 downto 0);
    signal type_cast_1312_wire : std_logic_vector(15 downto 0);
    signal type_cast_1316_wire : std_logic_vector(15 downto 0);
    signal type_cast_1318_wire : std_logic_vector(15 downto 0);
    signal type_cast_1323_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1325_wire : std_logic_vector(15 downto 0);
    signal type_cast_1332_wire : std_logic_vector(31 downto 0);
    signal type_cast_1336_wire : std_logic_vector(7 downto 0);
    signal type_cast_1345_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1385_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1390_wire : std_logic_vector(31 downto 0);
    signal type_cast_1393_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1400_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1405_wire : std_logic_vector(31 downto 0);
    signal type_cast_1408_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1424_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1429_wire : std_logic_vector(31 downto 0);
    signal type_cast_1432_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1439_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1445_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1455_wire : std_logic_vector(31 downto 0);
    signal type_cast_1458_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1467_wire : std_logic_vector(15 downto 0);
    signal type_cast_1469_wire : std_logic_vector(15 downto 0);
    signal type_cast_1474_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1476_wire : std_logic_vector(15 downto 0);
    signal type_cast_1481_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1483_wire : std_logic_vector(15 downto 0);
    signal type_cast_1487_wire : std_logic_vector(31 downto 0);
    signal type_cast_1492_wire : std_logic_vector(31 downto 0);
    signal type_cast_1494_wire : std_logic_vector(31 downto 0);
    signal type_cast_1514_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1524_wire : std_logic_vector(31 downto 0);
    signal type_cast_1526_wire : std_logic_vector(31 downto 0);
    signal type_cast_1538_wire : std_logic_vector(31 downto 0);
    signal type_cast_1543_wire : std_logic_vector(31 downto 0);
    signal type_cast_1545_wire : std_logic_vector(31 downto 0);
    signal type_cast_1569_wire : std_logic_vector(31 downto 0);
    signal type_cast_1571_wire : std_logic_vector(31 downto 0);
    signal type_cast_1583_wire : std_logic_vector(31 downto 0);
    signal type_cast_1588_wire : std_logic_vector(31 downto 0);
    signal type_cast_1613_wire : std_logic_vector(31 downto 0);
    signal type_cast_1616_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1622_wire : std_logic_vector(63 downto 0);
    signal type_cast_1635_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1641_wire : std_logic_vector(31 downto 0);
    signal type_cast_1696_wire : std_logic_vector(31 downto 0);
    signal type_cast_1699_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1705_wire : std_logic_vector(63 downto 0);
    signal type_cast_1721_wire : std_logic_vector(31 downto 0);
    signal type_cast_1724_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1730_wire : std_logic_vector(63 downto 0);
    signal type_cast_1748_wire : std_logic_vector(31 downto 0);
    signal type_cast_1754_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1759_wire : std_logic_vector(31 downto 0);
    signal type_cast_1761_wire : std_logic_vector(31 downto 0);
    signal type_cast_1774_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1782_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1787_wire : std_logic_vector(31 downto 0);
    signal type_cast_1824_wire : std_logic_vector(31 downto 0);
    signal type_cast_1837_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1860_wire : std_logic_vector(15 downto 0);
    signal type_cast_1862_wire : std_logic_vector(15 downto 0);
    signal type_cast_1866_wire : std_logic_vector(15 downto 0);
    signal type_cast_1868_wire : std_logic_vector(15 downto 0);
    signal type_cast_1872_wire : std_logic_vector(15 downto 0);
    signal type_cast_1875_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1882_wire : std_logic_vector(7 downto 0);
    signal type_cast_1886_wire : std_logic_vector(31 downto 0);
    signal type_cast_1895_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1935_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1940_wire : std_logic_vector(31 downto 0);
    signal type_cast_1943_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1950_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1955_wire : std_logic_vector(31 downto 0);
    signal type_cast_1958_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1974_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1979_wire : std_logic_vector(31 downto 0);
    signal type_cast_1982_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1989_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1995_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2005_wire : std_logic_vector(31 downto 0);
    signal type_cast_2008_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2017_wire : std_logic_vector(15 downto 0);
    signal type_cast_2020_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2024_wire : std_logic_vector(15 downto 0);
    signal type_cast_2026_wire : std_logic_vector(15 downto 0);
    signal type_cast_2030_wire : std_logic_vector(15 downto 0);
    signal type_cast_2033_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2037_wire : std_logic_vector(31 downto 0);
    signal type_cast_2042_wire : std_logic_vector(31 downto 0);
    signal type_cast_2044_wire : std_logic_vector(31 downto 0);
    signal type_cast_2064_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2074_wire : std_logic_vector(31 downto 0);
    signal type_cast_2076_wire : std_logic_vector(31 downto 0);
    signal type_cast_2088_wire : std_logic_vector(31 downto 0);
    signal type_cast_2093_wire : std_logic_vector(31 downto 0);
    signal type_cast_2095_wire : std_logic_vector(31 downto 0);
    signal type_cast_2115_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2125_wire : std_logic_vector(31 downto 0);
    signal type_cast_2127_wire : std_logic_vector(31 downto 0);
    signal type_cast_2139_wire : std_logic_vector(31 downto 0);
    signal type_cast_2144_wire : std_logic_vector(31 downto 0);
    signal type_cast_2169_wire : std_logic_vector(31 downto 0);
    signal type_cast_2172_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2178_wire : std_logic_vector(63 downto 0);
    signal type_cast_2191_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2197_wire : std_logic_vector(31 downto 0);
    signal type_cast_2252_wire : std_logic_vector(31 downto 0);
    signal type_cast_2255_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2261_wire : std_logic_vector(63 downto 0);
    signal type_cast_2277_wire : std_logic_vector(31 downto 0);
    signal type_cast_2280_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2286_wire : std_logic_vector(63 downto 0);
    signal type_cast_2304_wire : std_logic_vector(31 downto 0);
    signal type_cast_2310_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2315_wire : std_logic_vector(31 downto 0);
    signal type_cast_2317_wire : std_logic_vector(31 downto 0);
    signal type_cast_2330_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2338_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2343_wire : std_logic_vector(31 downto 0);
    signal type_cast_2356_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2381_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2387_wire : std_logic_vector(31 downto 0);
    signal type_cast_2400_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2423_wire : std_logic_vector(15 downto 0);
    signal type_cast_2426_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2430_wire : std_logic_vector(15 downto 0);
    signal type_cast_2432_wire : std_logic_vector(15 downto 0);
    signal type_cast_2436_wire : std_logic_vector(15 downto 0);
    signal type_cast_2438_wire : std_logic_vector(15 downto 0);
    signal type_cast_2445_wire : std_logic_vector(7 downto 0);
    signal type_cast_2449_wire : std_logic_vector(31 downto 0);
    signal type_cast_2453_wire : std_logic_vector(7 downto 0);
    signal type_cast_2462_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2472_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2512_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2517_wire : std_logic_vector(31 downto 0);
    signal type_cast_2520_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2527_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2532_wire : std_logic_vector(31 downto 0);
    signal type_cast_2535_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2551_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2556_wire : std_logic_vector(31 downto 0);
    signal type_cast_2559_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2566_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2572_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2582_wire : std_logic_vector(31 downto 0);
    signal type_cast_2585_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2595_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2597_wire : std_logic_vector(15 downto 0);
    signal type_cast_2601_wire : std_logic_vector(15 downto 0);
    signal type_cast_2603_wire : std_logic_vector(15 downto 0);
    signal type_cast_2607_wire : std_logic_vector(15 downto 0);
    signal type_cast_2609_wire : std_logic_vector(15 downto 0);
    signal type_cast_2613_wire : std_logic_vector(31 downto 0);
    signal type_cast_2618_wire : std_logic_vector(31 downto 0);
    signal type_cast_2620_wire : std_logic_vector(31 downto 0);
    signal type_cast_2640_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2650_wire : std_logic_vector(31 downto 0);
    signal type_cast_2652_wire : std_logic_vector(31 downto 0);
    signal type_cast_2664_wire : std_logic_vector(31 downto 0);
    signal type_cast_2669_wire : std_logic_vector(31 downto 0);
    signal type_cast_2671_wire : std_logic_vector(31 downto 0);
    signal type_cast_2695_wire : std_logic_vector(31 downto 0);
    signal type_cast_2697_wire : std_logic_vector(31 downto 0);
    signal type_cast_2709_wire : std_logic_vector(31 downto 0);
    signal type_cast_2714_wire : std_logic_vector(31 downto 0);
    signal type_cast_2739_wire : std_logic_vector(31 downto 0);
    signal type_cast_2742_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2748_wire : std_logic_vector(63 downto 0);
    signal type_cast_2761_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2767_wire : std_logic_vector(31 downto 0);
    signal type_cast_2822_wire : std_logic_vector(31 downto 0);
    signal type_cast_2825_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2831_wire : std_logic_vector(63 downto 0);
    signal type_cast_2847_wire : std_logic_vector(31 downto 0);
    signal type_cast_2850_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2856_wire : std_logic_vector(63 downto 0);
    signal type_cast_2874_wire : std_logic_vector(31 downto 0);
    signal type_cast_2880_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2885_wire : std_logic_vector(31 downto 0);
    signal type_cast_2887_wire : std_logic_vector(31 downto 0);
    signal type_cast_2900_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2908_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2913_wire : std_logic_vector(31 downto 0);
    signal type_cast_2950_wire : std_logic_vector(31 downto 0);
    signal type_cast_2963_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2986_wire : std_logic_vector(15 downto 0);
    signal type_cast_2989_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2993_wire : std_logic_vector(15 downto 0);
    signal type_cast_2995_wire : std_logic_vector(15 downto 0);
    signal type_cast_2999_wire : std_logic_vector(15 downto 0);
    signal type_cast_3001_wire : std_logic_vector(15 downto 0);
    signal type_cast_3008_wire : std_logic_vector(7 downto 0);
    signal type_cast_3012_wire : std_logic_vector(31 downto 0);
    signal type_cast_3021_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3061_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3066_wire : std_logic_vector(31 downto 0);
    signal type_cast_3069_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3076_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3081_wire : std_logic_vector(31 downto 0);
    signal type_cast_3084_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3100_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3105_wire : std_logic_vector(31 downto 0);
    signal type_cast_3108_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3115_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3121_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3131_wire : std_logic_vector(31 downto 0);
    signal type_cast_3134_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3144_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3146_wire : std_logic_vector(15 downto 0);
    signal type_cast_3150_wire : std_logic_vector(15 downto 0);
    signal type_cast_3152_wire : std_logic_vector(15 downto 0);
    signal type_cast_3156_wire : std_logic_vector(15 downto 0);
    signal type_cast_3159_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3163_wire : std_logic_vector(31 downto 0);
    signal type_cast_3168_wire : std_logic_vector(31 downto 0);
    signal type_cast_3170_wire : std_logic_vector(31 downto 0);
    signal type_cast_3190_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3196_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3206_wire : std_logic_vector(31 downto 0);
    signal type_cast_3208_wire : std_logic_vector(31 downto 0);
    signal type_cast_3220_wire : std_logic_vector(31 downto 0);
    signal type_cast_3225_wire : std_logic_vector(31 downto 0);
    signal type_cast_3227_wire : std_logic_vector(31 downto 0);
    signal type_cast_3247_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3257_wire : std_logic_vector(31 downto 0);
    signal type_cast_3259_wire : std_logic_vector(31 downto 0);
    signal type_cast_3271_wire : std_logic_vector(31 downto 0);
    signal type_cast_3276_wire : std_logic_vector(31 downto 0);
    signal type_cast_3301_wire : std_logic_vector(31 downto 0);
    signal type_cast_3304_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3310_wire : std_logic_vector(63 downto 0);
    signal type_cast_3323_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3329_wire : std_logic_vector(31 downto 0);
    signal type_cast_3384_wire : std_logic_vector(31 downto 0);
    signal type_cast_3387_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3393_wire : std_logic_vector(63 downto 0);
    signal type_cast_3409_wire : std_logic_vector(31 downto 0);
    signal type_cast_3412_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3418_wire : std_logic_vector(63 downto 0);
    signal type_cast_3436_wire : std_logic_vector(31 downto 0);
    signal type_cast_3442_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3447_wire : std_logic_vector(31 downto 0);
    signal type_cast_3449_wire : std_logic_vector(31 downto 0);
    signal type_cast_3462_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3470_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3475_wire : std_logic_vector(31 downto 0);
    signal type_cast_3488_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3513_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3519_wire : std_logic_vector(31 downto 0);
    signal type_cast_3532_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3538_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3561_wire : std_logic_vector(15 downto 0);
    signal type_cast_3564_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3568_wire : std_logic_vector(15 downto 0);
    signal type_cast_3570_wire : std_logic_vector(15 downto 0);
    signal type_cast_3574_wire : std_logic_vector(15 downto 0);
    signal type_cast_3576_wire : std_logic_vector(15 downto 0);
    signal type_cast_3583_wire : std_logic_vector(7 downto 0);
    signal type_cast_3587_wire : std_logic_vector(31 downto 0);
    signal type_cast_3591_wire : std_logic_vector(7 downto 0);
    signal type_cast_3600_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3610_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3650_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3655_wire : std_logic_vector(31 downto 0);
    signal type_cast_3658_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3665_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3670_wire : std_logic_vector(31 downto 0);
    signal type_cast_3673_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3689_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3694_wire : std_logic_vector(31 downto 0);
    signal type_cast_3697_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3704_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3710_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3720_wire : std_logic_vector(31 downto 0);
    signal type_cast_3723_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3732_wire : std_logic_vector(15 downto 0);
    signal type_cast_3735_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3739_wire : std_logic_vector(15 downto 0);
    signal type_cast_3741_wire : std_logic_vector(15 downto 0);
    signal type_cast_3745_wire : std_logic_vector(15 downto 0);
    signal type_cast_3747_wire : std_logic_vector(15 downto 0);
    signal type_cast_3751_wire : std_logic_vector(31 downto 0);
    signal type_cast_3756_wire : std_logic_vector(31 downto 0);
    signal type_cast_3758_wire : std_logic_vector(31 downto 0);
    signal type_cast_3778_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3784_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3794_wire : std_logic_vector(31 downto 0);
    signal type_cast_3796_wire : std_logic_vector(31 downto 0);
    signal type_cast_3808_wire : std_logic_vector(31 downto 0);
    signal type_cast_3813_wire : std_logic_vector(31 downto 0);
    signal type_cast_3815_wire : std_logic_vector(31 downto 0);
    signal type_cast_3839_wire : std_logic_vector(31 downto 0);
    signal type_cast_3841_wire : std_logic_vector(31 downto 0);
    signal type_cast_3853_wire : std_logic_vector(31 downto 0);
    signal type_cast_3858_wire : std_logic_vector(31 downto 0);
    signal type_cast_3883_wire : std_logic_vector(31 downto 0);
    signal type_cast_3886_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3892_wire : std_logic_vector(63 downto 0);
    signal type_cast_3905_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3911_wire : std_logic_vector(31 downto 0);
    signal type_cast_3966_wire : std_logic_vector(31 downto 0);
    signal type_cast_3969_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3975_wire : std_logic_vector(63 downto 0);
    signal type_cast_3991_wire : std_logic_vector(31 downto 0);
    signal type_cast_3994_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4000_wire : std_logic_vector(63 downto 0);
    signal type_cast_4018_wire : std_logic_vector(31 downto 0);
    signal type_cast_4024_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4029_wire : std_logic_vector(31 downto 0);
    signal type_cast_4031_wire : std_logic_vector(31 downto 0);
    signal type_cast_4044_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4052_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4057_wire : std_logic_vector(31 downto 0);
    signal type_cast_4094_wire : std_logic_vector(31 downto 0);
    signal type_cast_4107_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4113_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4136_wire : std_logic_vector(15 downto 0);
    signal type_cast_4139_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4143_wire : std_logic_vector(15 downto 0);
    signal type_cast_4145_wire : std_logic_vector(15 downto 0);
    signal type_cast_4149_wire : std_logic_vector(15 downto 0);
    signal type_cast_4151_wire : std_logic_vector(15 downto 0);
    signal type_cast_4158_wire : std_logic_vector(7 downto 0);
    signal type_cast_4162_wire : std_logic_vector(31 downto 0);
    signal type_cast_4171_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4177_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4217_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4222_wire : std_logic_vector(31 downto 0);
    signal type_cast_4225_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4232_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4237_wire : std_logic_vector(31 downto 0);
    signal type_cast_4240_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4256_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4261_wire : std_logic_vector(31 downto 0);
    signal type_cast_4264_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4271_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4277_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4287_wire : std_logic_vector(31 downto 0);
    signal type_cast_4290_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4300_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4302_wire : std_logic_vector(15 downto 0);
    signal type_cast_4306_wire : std_logic_vector(15 downto 0);
    signal type_cast_4308_wire : std_logic_vector(15 downto 0);
    signal type_cast_4313_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4315_wire : std_logic_vector(15 downto 0);
    signal type_cast_4319_wire : std_logic_vector(31 downto 0);
    signal type_cast_4324_wire : std_logic_vector(31 downto 0);
    signal type_cast_4326_wire : std_logic_vector(31 downto 0);
    signal type_cast_4350_wire : std_logic_vector(31 downto 0);
    signal type_cast_4352_wire : std_logic_vector(31 downto 0);
    signal type_cast_4364_wire : std_logic_vector(31 downto 0);
    signal type_cast_4369_wire : std_logic_vector(31 downto 0);
    signal type_cast_4371_wire : std_logic_vector(31 downto 0);
    signal type_cast_4391_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4401_wire : std_logic_vector(31 downto 0);
    signal type_cast_4403_wire : std_logic_vector(31 downto 0);
    signal type_cast_4415_wire : std_logic_vector(31 downto 0);
    signal type_cast_4420_wire : std_logic_vector(31 downto 0);
    signal type_cast_4445_wire : std_logic_vector(31 downto 0);
    signal type_cast_4448_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4454_wire : std_logic_vector(63 downto 0);
    signal type_cast_4467_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_4473_wire : std_logic_vector(31 downto 0);
    signal type_cast_4528_wire : std_logic_vector(31 downto 0);
    signal type_cast_4531_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4537_wire : std_logic_vector(63 downto 0);
    signal type_cast_4553_wire : std_logic_vector(31 downto 0);
    signal type_cast_4556_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4562_wire : std_logic_vector(63 downto 0);
    signal type_cast_4580_wire : std_logic_vector(31 downto 0);
    signal type_cast_4586_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4591_wire : std_logic_vector(31 downto 0);
    signal type_cast_4593_wire : std_logic_vector(31 downto 0);
    signal type_cast_4606_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4614_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4619_wire : std_logic_vector(31 downto 0);
    signal type_cast_4632_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4657_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4663_wire : std_logic_vector(31 downto 0);
    signal type_cast_4694_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4696_wire : std_logic_vector(15 downto 0);
    signal type_cast_4700_wire : std_logic_vector(15 downto 0);
    signal type_cast_4702_wire : std_logic_vector(15 downto 0);
    signal type_cast_4706_wire : std_logic_vector(15 downto 0);
    signal type_cast_4708_wire : std_logic_vector(15 downto 0);
    signal type_cast_4715_wire : std_logic_vector(7 downto 0);
    signal type_cast_4719_wire : std_logic_vector(31 downto 0);
    signal type_cast_4723_wire : std_logic_vector(7 downto 0);
    signal type_cast_4732_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4742_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4748_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4788_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4793_wire : std_logic_vector(31 downto 0);
    signal type_cast_4796_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4803_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4808_wire : std_logic_vector(31 downto 0);
    signal type_cast_4811_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4827_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4832_wire : std_logic_vector(31 downto 0);
    signal type_cast_4835_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4842_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4848_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4858_wire : std_logic_vector(31 downto 0);
    signal type_cast_4861_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4871_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4873_wire : std_logic_vector(15 downto 0);
    signal type_cast_4877_wire : std_logic_vector(15 downto 0);
    signal type_cast_4879_wire : std_logic_vector(15 downto 0);
    signal type_cast_4883_wire : std_logic_vector(15 downto 0);
    signal type_cast_4885_wire : std_logic_vector(15 downto 0);
    signal type_cast_4889_wire : std_logic_vector(31 downto 0);
    signal type_cast_4894_wire : std_logic_vector(31 downto 0);
    signal type_cast_4896_wire : std_logic_vector(31 downto 0);
    signal type_cast_4920_wire : std_logic_vector(31 downto 0);
    signal type_cast_4922_wire : std_logic_vector(31 downto 0);
    signal type_cast_4934_wire : std_logic_vector(31 downto 0);
    signal type_cast_4939_wire : std_logic_vector(31 downto 0);
    signal type_cast_4941_wire : std_logic_vector(31 downto 0);
    signal type_cast_4965_wire : std_logic_vector(31 downto 0);
    signal type_cast_4967_wire : std_logic_vector(31 downto 0);
    signal type_cast_4979_wire : std_logic_vector(31 downto 0);
    signal type_cast_4984_wire : std_logic_vector(31 downto 0);
    signal type_cast_5009_wire : std_logic_vector(31 downto 0);
    signal type_cast_5012_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_5018_wire : std_logic_vector(63 downto 0);
    signal type_cast_5031_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_5037_wire : std_logic_vector(31 downto 0);
    signal type_cast_5092_wire : std_logic_vector(31 downto 0);
    signal type_cast_5095_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_5101_wire : std_logic_vector(63 downto 0);
    signal type_cast_5117_wire : std_logic_vector(31 downto 0);
    signal type_cast_5120_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_5126_wire : std_logic_vector(63 downto 0);
    signal type_cast_5144_wire : std_logic_vector(31 downto 0);
    signal type_cast_5150_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_5155_wire : std_logic_vector(31 downto 0);
    signal type_cast_5157_wire : std_logic_vector(31 downto 0);
    signal type_cast_5170_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_5178_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_5183_wire : std_logic_vector(31 downto 0);
    signal type_cast_5220_wire : std_logic_vector(31 downto 0);
    signal type_cast_5250_wire : std_logic_vector(15 downto 0);
    signal type_cast_5253_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_5257_wire : std_logic_vector(15 downto 0);
    signal type_cast_5259_wire : std_logic_vector(15 downto 0);
    signal type_cast_5263_wire : std_logic_vector(15 downto 0);
    signal type_cast_5265_wire : std_logic_vector(15 downto 0);
    signal type_cast_819_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_825_wire : std_logic_vector(31 downto 0);
    signal type_cast_828_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_835_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_840_wire : std_logic_vector(31 downto 0);
    signal type_cast_843_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_859_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_864_wire : std_logic_vector(31 downto 0);
    signal type_cast_867_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_874_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_880_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_890_wire : std_logic_vector(31 downto 0);
    signal type_cast_893_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_903_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_905_wire : std_logic_vector(15 downto 0);
    signal type_cast_910_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_912_wire : std_logic_vector(15 downto 0);
    signal type_cast_917_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_919_wire : std_logic_vector(15 downto 0);
    signal type_cast_923_wire : std_logic_vector(31 downto 0);
    signal type_cast_928_wire : std_logic_vector(31 downto 0);
    signal type_cast_930_wire : std_logic_vector(31 downto 0);
    signal type_cast_950_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_960_wire : std_logic_vector(31 downto 0);
    signal type_cast_962_wire : std_logic_vector(31 downto 0);
    signal type_cast_974_wire : std_logic_vector(31 downto 0);
    signal type_cast_979_wire : std_logic_vector(31 downto 0);
    signal type_cast_981_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_col_high_1234_word_address_0 <= "0";
    LOAD_col_high_1556_word_address_0 <= "0";
    LOAD_col_high_1791_word_address_0 <= "0";
    LOAD_col_high_2106_word_address_0 <= "0";
    LOAD_col_high_2347_word_address_0 <= "0";
    LOAD_col_high_2682_word_address_0 <= "0";
    LOAD_col_high_2917_word_address_0 <= "0";
    LOAD_col_high_3238_word_address_0 <= "0";
    LOAD_col_high_3479_word_address_0 <= "0";
    LOAD_col_high_3826_word_address_0 <= "0";
    LOAD_col_high_4061_word_address_0 <= "0";
    LOAD_col_high_4382_word_address_0 <= "0";
    LOAD_col_high_4623_word_address_0 <= "0";
    LOAD_col_high_4952_word_address_0 <= "0";
    LOAD_col_high_5187_word_address_0 <= "0";
    LOAD_col_high_782_word_address_0 <= "0";
    LOAD_col_high_992_word_address_0 <= "0";
    LOAD_depth_high_1352_word_address_0 <= "0";
    LOAD_depth_high_1902_word_address_0 <= "0";
    LOAD_depth_high_2479_word_address_0 <= "0";
    LOAD_depth_high_3028_word_address_0 <= "0";
    LOAD_depth_high_3617_word_address_0 <= "0";
    LOAD_depth_high_4184_word_address_0 <= "0";
    LOAD_depth_high_4755_word_address_0 <= "0";
    LOAD_depth_high_779_word_address_0 <= "0";
    LOAD_pad_1349_word_address_0 <= "0";
    LOAD_pad_1899_word_address_0 <= "0";
    LOAD_pad_2476_word_address_0 <= "0";
    LOAD_pad_3025_word_address_0 <= "0";
    LOAD_pad_3614_word_address_0 <= "0";
    LOAD_pad_4181_word_address_0 <= "0";
    LOAD_pad_4752_word_address_0 <= "0";
    LOAD_pad_776_word_address_0 <= "0";
    LOAD_row_high_1278_word_address_0 <= "0";
    LOAD_row_high_1505_word_address_0 <= "0";
    LOAD_row_high_1828_word_address_0 <= "0";
    LOAD_row_high_2055_word_address_0 <= "0";
    LOAD_row_high_2391_word_address_0 <= "0";
    LOAD_row_high_2631_word_address_0 <= "0";
    LOAD_row_high_2954_word_address_0 <= "0";
    LOAD_row_high_3181_word_address_0 <= "0";
    LOAD_row_high_3523_word_address_0 <= "0";
    LOAD_row_high_3769_word_address_0 <= "0";
    LOAD_row_high_4098_word_address_0 <= "0";
    LOAD_row_high_4337_word_address_0 <= "0";
    LOAD_row_high_4667_word_address_0 <= "0";
    LOAD_row_high_4907_word_address_0 <= "0";
    LOAD_row_high_5224_word_address_0 <= "0";
    LOAD_row_high_941_word_address_0 <= "0";
    STORE_col_high_752_word_address_0 <= "0";
    STORE_depth_high_771_word_address_0 <= "0";
    STORE_row_high_733_word_address_0 <= "0";
    array_obj_ref_1072_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1072_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1072_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1072_resized_base_address <= "00000000000000";
    array_obj_ref_1155_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1155_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1155_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1155_resized_base_address <= "00000000000000";
    array_obj_ref_1180_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1180_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1180_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1180_resized_base_address <= "00000000000000";
    array_obj_ref_1629_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1629_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1629_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1629_resized_base_address <= "00000000000000";
    array_obj_ref_1712_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1712_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1712_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1712_resized_base_address <= "00000000000000";
    array_obj_ref_1737_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1737_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1737_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1737_resized_base_address <= "00000000000000";
    array_obj_ref_2185_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2185_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2185_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2185_resized_base_address <= "00000000000000";
    array_obj_ref_2268_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2268_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2268_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2268_resized_base_address <= "00000000000000";
    array_obj_ref_2293_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2293_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2293_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2293_resized_base_address <= "00000000000000";
    array_obj_ref_2755_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2755_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2755_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2755_resized_base_address <= "00000000000000";
    array_obj_ref_2838_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2838_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2838_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2838_resized_base_address <= "00000000000000";
    array_obj_ref_2863_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2863_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2863_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2863_resized_base_address <= "00000000000000";
    array_obj_ref_3317_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3317_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3317_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3317_resized_base_address <= "00000000000000";
    array_obj_ref_3400_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3400_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3400_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3400_resized_base_address <= "00000000000000";
    array_obj_ref_3425_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3425_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3425_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3425_resized_base_address <= "00000000000000";
    array_obj_ref_3899_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3899_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3899_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3899_resized_base_address <= "00000000000000";
    array_obj_ref_3982_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3982_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3982_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3982_resized_base_address <= "00000000000000";
    array_obj_ref_4007_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4007_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4007_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4007_resized_base_address <= "00000000000000";
    array_obj_ref_4461_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4461_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4461_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4461_resized_base_address <= "00000000000000";
    array_obj_ref_4544_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4544_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4544_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4544_resized_base_address <= "00000000000000";
    array_obj_ref_4569_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4569_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4569_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4569_resized_base_address <= "00000000000000";
    array_obj_ref_5025_constant_part_of_offset <= "00000000000000";
    array_obj_ref_5025_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_5025_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_5025_resized_base_address <= "00000000000000";
    array_obj_ref_5108_constant_part_of_offset <= "00000000000000";
    array_obj_ref_5108_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_5108_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_5108_resized_base_address <= "00000000000000";
    array_obj_ref_5133_constant_part_of_offset <= "00000000000000";
    array_obj_ref_5133_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_5133_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_5133_resized_base_address <= "00000000000000";
    iNsTr_0_724 <= "00000000000000000000000000000011";
    iNsTr_101_4193 <= "00000000000000000000000000000101";
    iNsTr_102_4205 <= "00000000000000000000000000000100";
    iNsTr_117_4764 <= "00000000000000000000000000000101";
    iNsTr_118_4776 <= "00000000000000000000000000000100";
    iNsTr_21_1361 <= "00000000000000000000000000000101";
    iNsTr_22_1373 <= "00000000000000000000000000000100";
    iNsTr_2_743 <= "00000000000000000000000000000100";
    iNsTr_37_1911 <= "00000000000000000000000000000101";
    iNsTr_38_1923 <= "00000000000000000000000000000100";
    iNsTr_4_762 <= "00000000000000000000000000000101";
    iNsTr_53_2488 <= "00000000000000000000000000000101";
    iNsTr_54_2500 <= "00000000000000000000000000000100";
    iNsTr_69_3037 <= "00000000000000000000000000000101";
    iNsTr_70_3049 <= "00000000000000000000000000000100";
    iNsTr_7_791 <= "00000000000000000000000000000101";
    iNsTr_85_3626 <= "00000000000000000000000000000101";
    iNsTr_86_3638 <= "00000000000000000000000000000100";
    iNsTr_8_803 <= "00000000000000000000000000000100";
    ptr_deref_1076_word_offset_0 <= "00000000000000";
    ptr_deref_1160_word_offset_0 <= "00000000000000";
    ptr_deref_1184_word_offset_0 <= "00000000000000";
    ptr_deref_1364_word_offset_0 <= "0000000";
    ptr_deref_1376_word_offset_0 <= "0000000";
    ptr_deref_1633_word_offset_0 <= "00000000000000";
    ptr_deref_1717_word_offset_0 <= "00000000000000";
    ptr_deref_1741_word_offset_0 <= "00000000000000";
    ptr_deref_1914_word_offset_0 <= "0000000";
    ptr_deref_1926_word_offset_0 <= "0000000";
    ptr_deref_2189_word_offset_0 <= "00000000000000";
    ptr_deref_2273_word_offset_0 <= "00000000000000";
    ptr_deref_2297_word_offset_0 <= "00000000000000";
    ptr_deref_2491_word_offset_0 <= "0000000";
    ptr_deref_2503_word_offset_0 <= "0000000";
    ptr_deref_2759_word_offset_0 <= "00000000000000";
    ptr_deref_2843_word_offset_0 <= "00000000000000";
    ptr_deref_2867_word_offset_0 <= "00000000000000";
    ptr_deref_3040_word_offset_0 <= "0000000";
    ptr_deref_3052_word_offset_0 <= "0000000";
    ptr_deref_3321_word_offset_0 <= "00000000000000";
    ptr_deref_3405_word_offset_0 <= "00000000000000";
    ptr_deref_3429_word_offset_0 <= "00000000000000";
    ptr_deref_3629_word_offset_0 <= "0000000";
    ptr_deref_3641_word_offset_0 <= "0000000";
    ptr_deref_3903_word_offset_0 <= "00000000000000";
    ptr_deref_3987_word_offset_0 <= "00000000000000";
    ptr_deref_4011_word_offset_0 <= "00000000000000";
    ptr_deref_4196_word_offset_0 <= "0000000";
    ptr_deref_4208_word_offset_0 <= "0000000";
    ptr_deref_4465_word_offset_0 <= "00000000000000";
    ptr_deref_4549_word_offset_0 <= "00000000000000";
    ptr_deref_4573_word_offset_0 <= "00000000000000";
    ptr_deref_4767_word_offset_0 <= "0000000";
    ptr_deref_4779_word_offset_0 <= "0000000";
    ptr_deref_5029_word_offset_0 <= "00000000000000";
    ptr_deref_5113_word_offset_0 <= "00000000000000";
    ptr_deref_5137_word_offset_0 <= "00000000000000";
    ptr_deref_727_word_offset_0 <= "0000000";
    ptr_deref_746_word_offset_0 <= "0000000";
    ptr_deref_765_word_offset_0 <= "0000000";
    ptr_deref_794_word_offset_0 <= "0000000";
    ptr_deref_806_word_offset_0 <= "0000000";
    type_cast_1001_wire_constant <= "00000000000000000000000000000001";
    type_cast_1058_wire_constant <= "00000000000000000000000000000010";
    type_cast_1078_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1142_wire_constant <= "00000000000000000000000000000010";
    type_cast_1167_wire_constant <= "00000000000000000000000000000010";
    type_cast_1197_wire_constant <= "00000000000000000000000000000100";
    type_cast_1217_wire_constant <= "0000000000000100";
    type_cast_1225_wire_constant <= "0000000000000001";
    type_cast_1243_wire_constant <= "00000000000000000000000000000001";
    type_cast_1268_wire_constant <= "0000000000000000";
    type_cast_1287_wire_constant <= "00000000000000000000000000000010";
    type_cast_1323_wire_constant <= "0000000000000000";
    type_cast_1345_wire_constant <= "0000000000000001";
    type_cast_1385_wire_constant <= "00000000000000000000000000010000";
    type_cast_1393_wire_constant <= "00000000000000000000000000010000";
    type_cast_1400_wire_constant <= "00000000000000000000000000010000";
    type_cast_1408_wire_constant <= "00000000000000000000000000010000";
    type_cast_1424_wire_constant <= "00000000000000000000000000010000";
    type_cast_1432_wire_constant <= "00000000000000000000000000010000";
    type_cast_1439_wire_constant <= "00000000000000000000000000000001";
    type_cast_1445_wire_constant <= "00000000000000000000000000010000";
    type_cast_1458_wire_constant <= "00000000000000000000000000010000";
    type_cast_1474_wire_constant <= "0000000000000000";
    type_cast_1481_wire_constant <= "0000000000000000";
    type_cast_1514_wire_constant <= "00000000000000000000000000000010";
    type_cast_1616_wire_constant <= "00000000000000000000000000000010";
    type_cast_1635_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1699_wire_constant <= "00000000000000000000000000000010";
    type_cast_1724_wire_constant <= "00000000000000000000000000000010";
    type_cast_1754_wire_constant <= "00000000000000000000000000000100";
    type_cast_1774_wire_constant <= "0000000000000100";
    type_cast_1782_wire_constant <= "0000000000000001";
    type_cast_1837_wire_constant <= "00000000000000000000000000000010";
    type_cast_1875_wire_constant <= "0000000000000000";
    type_cast_1895_wire_constant <= "0000000000000010";
    type_cast_1935_wire_constant <= "00000000000000000000000000010000";
    type_cast_1943_wire_constant <= "00000000000000000000000000010000";
    type_cast_1950_wire_constant <= "00000000000000000000000000010000";
    type_cast_1958_wire_constant <= "00000000000000000000000000010000";
    type_cast_1974_wire_constant <= "00000000000000000000000000010000";
    type_cast_1982_wire_constant <= "00000000000000000000000000010000";
    type_cast_1989_wire_constant <= "00000000000000000000000000000001";
    type_cast_1995_wire_constant <= "00000000000000000000000000010000";
    type_cast_2008_wire_constant <= "00000000000000000000000000010000";
    type_cast_2020_wire_constant <= "0000000000000000";
    type_cast_2033_wire_constant <= "0000000000000000";
    type_cast_2064_wire_constant <= "00000000000000000000000000000001";
    type_cast_2115_wire_constant <= "00000000000000000000000000000001";
    type_cast_2172_wire_constant <= "00000000000000000000000000000010";
    type_cast_2191_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2255_wire_constant <= "00000000000000000000000000000010";
    type_cast_2280_wire_constant <= "00000000000000000000000000000010";
    type_cast_2310_wire_constant <= "00000000000000000000000000000100";
    type_cast_2330_wire_constant <= "0000000000000100";
    type_cast_2338_wire_constant <= "0000000000000001";
    type_cast_2356_wire_constant <= "00000000000000000000000000000001";
    type_cast_2381_wire_constant <= "0000000000000000";
    type_cast_2400_wire_constant <= "00000000000000000000000000000001";
    type_cast_2426_wire_constant <= "0000000000000000";
    type_cast_2462_wire_constant <= "0000000000000001";
    type_cast_2472_wire_constant <= "0000000000000010";
    type_cast_2512_wire_constant <= "00000000000000000000000000010000";
    type_cast_2520_wire_constant <= "00000000000000000000000000010000";
    type_cast_2527_wire_constant <= "00000000000000000000000000010000";
    type_cast_2535_wire_constant <= "00000000000000000000000000010000";
    type_cast_2551_wire_constant <= "00000000000000000000000000010000";
    type_cast_2559_wire_constant <= "00000000000000000000000000010000";
    type_cast_2566_wire_constant <= "00000000000000000000000000000001";
    type_cast_2572_wire_constant <= "00000000000000000000000000010000";
    type_cast_2585_wire_constant <= "00000000000000000000000000010000";
    type_cast_2595_wire_constant <= "0000000000000000";
    type_cast_2640_wire_constant <= "00000000000000000000000000000001";
    type_cast_2742_wire_constant <= "00000000000000000000000000000010";
    type_cast_2761_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2825_wire_constant <= "00000000000000000000000000000010";
    type_cast_2850_wire_constant <= "00000000000000000000000000000010";
    type_cast_2880_wire_constant <= "00000000000000000000000000000100";
    type_cast_2900_wire_constant <= "0000000000000100";
    type_cast_2908_wire_constant <= "0000000000000001";
    type_cast_2963_wire_constant <= "00000000000000000000000000000001";
    type_cast_2989_wire_constant <= "0000000000000000";
    type_cast_3021_wire_constant <= "0000000000000001";
    type_cast_3061_wire_constant <= "00000000000000000000000000010000";
    type_cast_3069_wire_constant <= "00000000000000000000000000010000";
    type_cast_3076_wire_constant <= "00000000000000000000000000010000";
    type_cast_3084_wire_constant <= "00000000000000000000000000010000";
    type_cast_3100_wire_constant <= "00000000000000000000000000010000";
    type_cast_3108_wire_constant <= "00000000000000000000000000010000";
    type_cast_3115_wire_constant <= "00000000000000000000000000000001";
    type_cast_3121_wire_constant <= "00000000000000000000000000010000";
    type_cast_3134_wire_constant <= "00000000000000000000000000010000";
    type_cast_3144_wire_constant <= "0000000000000000";
    type_cast_3159_wire_constant <= "0000000000000000";
    type_cast_3190_wire_constant <= "00000000000000000000000000000011";
    type_cast_3196_wire_constant <= "00000000000000000000000000000010";
    type_cast_3247_wire_constant <= "00000000000000000000000000000001";
    type_cast_3304_wire_constant <= "00000000000000000000000000000010";
    type_cast_3323_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_3387_wire_constant <= "00000000000000000000000000000010";
    type_cast_3412_wire_constant <= "00000000000000000000000000000010";
    type_cast_3442_wire_constant <= "00000000000000000000000000000100";
    type_cast_3462_wire_constant <= "0000000000000100";
    type_cast_3470_wire_constant <= "0000000000000001";
    type_cast_3488_wire_constant <= "00000000000000000000000000000001";
    type_cast_3513_wire_constant <= "0000000000000000";
    type_cast_3532_wire_constant <= "00000000000000000000000000000011";
    type_cast_3538_wire_constant <= "00000000000000000000000000000010";
    type_cast_3564_wire_constant <= "0000000000000000";
    type_cast_3600_wire_constant <= "0000000000000001";
    type_cast_3610_wire_constant <= "0000000000000001";
    type_cast_3650_wire_constant <= "00000000000000000000000000010000";
    type_cast_3658_wire_constant <= "00000000000000000000000000010000";
    type_cast_3665_wire_constant <= "00000000000000000000000000010000";
    type_cast_3673_wire_constant <= "00000000000000000000000000010000";
    type_cast_3689_wire_constant <= "00000000000000000000000000010000";
    type_cast_3697_wire_constant <= "00000000000000000000000000010000";
    type_cast_3704_wire_constant <= "00000000000000000000000000000001";
    type_cast_3710_wire_constant <= "00000000000000000000000000010000";
    type_cast_3723_wire_constant <= "00000000000000000000000000010000";
    type_cast_3735_wire_constant <= "0000000000000000";
    type_cast_3778_wire_constant <= "00000000000000000000000000000011";
    type_cast_3784_wire_constant <= "00000000000000000000000000000010";
    type_cast_3886_wire_constant <= "00000000000000000000000000000010";
    type_cast_3905_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_3969_wire_constant <= "00000000000000000000000000000010";
    type_cast_3994_wire_constant <= "00000000000000000000000000000010";
    type_cast_4024_wire_constant <= "00000000000000000000000000000100";
    type_cast_4044_wire_constant <= "0000000000000100";
    type_cast_4052_wire_constant <= "0000000000000001";
    type_cast_4107_wire_constant <= "00000000000000000000000000000011";
    type_cast_4113_wire_constant <= "00000000000000000000000000000010";
    type_cast_4139_wire_constant <= "0000000000000000";
    type_cast_4171_wire_constant <= "0000000000000010";
    type_cast_4177_wire_constant <= "0000000000000011";
    type_cast_4217_wire_constant <= "00000000000000000000000000010000";
    type_cast_4225_wire_constant <= "00000000000000000000000000010000";
    type_cast_4232_wire_constant <= "00000000000000000000000000010000";
    type_cast_4240_wire_constant <= "00000000000000000000000000010000";
    type_cast_4256_wire_constant <= "00000000000000000000000000010000";
    type_cast_4264_wire_constant <= "00000000000000000000000000010000";
    type_cast_4271_wire_constant <= "00000000000000000000000000000001";
    type_cast_4277_wire_constant <= "00000000000000000000000000010000";
    type_cast_4290_wire_constant <= "00000000000000000000000000010000";
    type_cast_4300_wire_constant <= "0000000000000000";
    type_cast_4313_wire_constant <= "0000000000000000";
    type_cast_4391_wire_constant <= "00000000000000000000000000000001";
    type_cast_4448_wire_constant <= "00000000000000000000000000000010";
    type_cast_4467_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_4531_wire_constant <= "00000000000000000000000000000010";
    type_cast_4556_wire_constant <= "00000000000000000000000000000010";
    type_cast_4586_wire_constant <= "00000000000000000000000000000100";
    type_cast_4606_wire_constant <= "0000000000000100";
    type_cast_4614_wire_constant <= "0000000000000001";
    type_cast_4632_wire_constant <= "00000000000000000000000000000001";
    type_cast_4657_wire_constant <= "0000000000000000";
    type_cast_4694_wire_constant <= "0000000000000000";
    type_cast_4732_wire_constant <= "0000000000000001";
    type_cast_4742_wire_constant <= "0000000000000011";
    type_cast_4748_wire_constant <= "0000000000000010";
    type_cast_4788_wire_constant <= "00000000000000000000000000010000";
    type_cast_4796_wire_constant <= "00000000000000000000000000010000";
    type_cast_4803_wire_constant <= "00000000000000000000000000010000";
    type_cast_4811_wire_constant <= "00000000000000000000000000010000";
    type_cast_4827_wire_constant <= "00000000000000000000000000010000";
    type_cast_4835_wire_constant <= "00000000000000000000000000010000";
    type_cast_4842_wire_constant <= "00000000000000000000000000000001";
    type_cast_4848_wire_constant <= "00000000000000000000000000010000";
    type_cast_4861_wire_constant <= "00000000000000000000000000010000";
    type_cast_4871_wire_constant <= "0000000000000000";
    type_cast_5012_wire_constant <= "00000000000000000000000000000010";
    type_cast_5031_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_5095_wire_constant <= "00000000000000000000000000000010";
    type_cast_5120_wire_constant <= "00000000000000000000000000000010";
    type_cast_5150_wire_constant <= "00000000000000000000000000000100";
    type_cast_5170_wire_constant <= "0000000000000100";
    type_cast_5178_wire_constant <= "0000000000000001";
    type_cast_5253_wire_constant <= "0000000000000000";
    type_cast_819_wire_constant <= "00000000000000000000000000010000";
    type_cast_828_wire_constant <= "00000000000000000000000000010000";
    type_cast_835_wire_constant <= "00000000000000000000000000010000";
    type_cast_843_wire_constant <= "00000000000000000000000000010000";
    type_cast_859_wire_constant <= "00000000000000000000000000010000";
    type_cast_867_wire_constant <= "00000000000000000000000000010000";
    type_cast_874_wire_constant <= "00000000000000000000000000000001";
    type_cast_880_wire_constant <= "00000000000000000000000000010000";
    type_cast_893_wire_constant <= "00000000000000000000000000010000";
    type_cast_903_wire_constant <= "0000000000000000";
    type_cast_910_wire_constant <= "0000000000000000";
    type_cast_917_wire_constant <= "0000000000000000";
    type_cast_950_wire_constant <= "00000000000000000000000000000010";
    phi_stmt_1307: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1310_wire & type_cast_1312_wire;
      req <= phi_stmt_1307_req_0 & phi_stmt_1307_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1307",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1307_ack_0,
          idata => idata,
          odata => jx_x0x_xph_1307,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1307
    phi_stmt_1313: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1316_wire & type_cast_1318_wire;
      req <= phi_stmt_1313_req_0 & phi_stmt_1313_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1313",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1313_ack_0,
          idata => idata,
          odata => ix_x1x_xph_1313,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1313
    phi_stmt_1319: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1323_wire_constant & type_cast_1325_wire;
      req <= phi_stmt_1319_req_0 & phi_stmt_1319_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1319",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1319_ack_0,
          idata => idata,
          odata => kx_x0x_xph_1319,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1319
    phi_stmt_1329: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1332_wire;
      req(0) <= phi_stmt_1329_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1329",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1329_ack_0,
          idata => idata,
          odata => conv155x_xlcssa_1329,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1329
    phi_stmt_1333: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1336_wire;
      req(0) <= phi_stmt_1333_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1333",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1333_ack_0,
          idata => idata,
          odata => tmp154x_xlcssa_1333,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1333
    phi_stmt_1464: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1467_wire & type_cast_1469_wire;
      req <= phi_stmt_1464_req_0 & phi_stmt_1464_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1464",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1464_ack_0,
          idata => idata,
          odata => j240x_x1_1464,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1464
    phi_stmt_1470: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1474_wire_constant & type_cast_1476_wire;
      req <= phi_stmt_1470_req_0 & phi_stmt_1470_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1470",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1470_ack_0,
          idata => idata,
          odata => i194x_x2_1470,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1470
    phi_stmt_1477: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1481_wire_constant & type_cast_1483_wire;
      req <= phi_stmt_1477_req_0 & phi_stmt_1477_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1477",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1477_ack_0,
          idata => idata,
          odata => k186x_x1_1477,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1477
    phi_stmt_1857: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1860_wire & type_cast_1862_wire;
      req <= phi_stmt_1857_req_0 & phi_stmt_1857_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1857",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1857_ack_0,
          idata => idata,
          odata => j240x_x0x_xph_1857,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1857
    phi_stmt_1863: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1866_wire & type_cast_1868_wire;
      req <= phi_stmt_1863_req_0 & phi_stmt_1863_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1863",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1863_ack_0,
          idata => idata,
          odata => i194x_x1x_xph_1863,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1863
    phi_stmt_1869: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1872_wire & type_cast_1875_wire_constant;
      req <= phi_stmt_1869_req_0 & phi_stmt_1869_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1869",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1869_ack_0,
          idata => idata,
          odata => k186x_x0x_xph_1869,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1869
    phi_stmt_1879: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1882_wire;
      req(0) <= phi_stmt_1879_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1879",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1879_ack_0,
          idata => idata,
          odata => tmp383x_xlcssa_1879,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1879
    phi_stmt_1883: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1886_wire;
      req(0) <= phi_stmt_1883_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1883",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1883_ack_0,
          idata => idata,
          odata => conv369x_xlcssa_1883,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1883
    phi_stmt_2014: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2017_wire & type_cast_2020_wire_constant;
      req <= phi_stmt_2014_req_0 & phi_stmt_2014_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2014",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2014_ack_0,
          idata => idata,
          odata => k402x_x1_2014,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2014
    phi_stmt_2021: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2024_wire & type_cast_2026_wire;
      req <= phi_stmt_2021_req_0 & phi_stmt_2021_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2021",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2021_ack_0,
          idata => idata,
          odata => i406x_x2_2021,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2021
    phi_stmt_2027: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2030_wire & type_cast_2033_wire_constant;
      req <= phi_stmt_2027_req_0 & phi_stmt_2027_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2027",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2027_ack_0,
          idata => idata,
          odata => j456x_x1_2027,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2027
    phi_stmt_2420: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2423_wire & type_cast_2426_wire_constant;
      req <= phi_stmt_2420_req_0 & phi_stmt_2420_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2420",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2420_ack_0,
          idata => idata,
          odata => k402x_x0x_xph_2420,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2420
    phi_stmt_2427: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2430_wire & type_cast_2432_wire;
      req <= phi_stmt_2427_req_0 & phi_stmt_2427_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2427",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2427_ack_0,
          idata => idata,
          odata => i406x_x1x_xph_2427,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2427
    phi_stmt_2433: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2436_wire & type_cast_2438_wire;
      req <= phi_stmt_2433_req_0 & phi_stmt_2433_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2433",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2433_ack_0,
          idata => idata,
          odata => j456x_x0x_xph_2433,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2433
    phi_stmt_2442: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2445_wire;
      req(0) <= phi_stmt_2442_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2442",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2442_ack_0,
          idata => idata,
          odata => tmp601x_xlcssa_2442,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2442
    phi_stmt_2446: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2449_wire;
      req(0) <= phi_stmt_2446_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2446",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2446_ack_0,
          idata => idata,
          odata => conv586x_xlcssa_2446,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2446
    phi_stmt_2450: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2453_wire;
      req(0) <= phi_stmt_2450_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2450",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2450_ack_0,
          idata => idata,
          odata => tmp585x_xlcssa_2450,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2450
    phi_stmt_2591: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2595_wire_constant & type_cast_2597_wire;
      req <= phi_stmt_2591_req_0 & phi_stmt_2591_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2591",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2591_ack_0,
          idata => idata,
          odata => k620x_x1_2591,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2591
    phi_stmt_2598: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2601_wire & type_cast_2603_wire;
      req <= phi_stmt_2598_req_0 & phi_stmt_2598_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2598",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2598_ack_0,
          idata => idata,
          odata => i628x_x2_2598,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2598
    phi_stmt_2604: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2607_wire & type_cast_2609_wire;
      req <= phi_stmt_2604_req_0 & phi_stmt_2604_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2604",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2604_ack_0,
          idata => idata,
          odata => j678x_x1_2604,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2604
    phi_stmt_2983: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2986_wire & type_cast_2989_wire_constant;
      req <= phi_stmt_2983_req_0 & phi_stmt_2983_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2983",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2983_ack_0,
          idata => idata,
          odata => k620x_x0x_xph_2983,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2983
    phi_stmt_2990: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2993_wire & type_cast_2995_wire;
      req <= phi_stmt_2990_req_0 & phi_stmt_2990_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2990",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2990_ack_0,
          idata => idata,
          odata => i628x_x1x_xph_2990,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2990
    phi_stmt_2996: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2999_wire & type_cast_3001_wire;
      req <= phi_stmt_2996_req_0 & phi_stmt_2996_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2996",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2996_ack_0,
          idata => idata,
          odata => j678x_x0x_xph_2996,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2996
    phi_stmt_3005: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3008_wire;
      req(0) <= phi_stmt_3005_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3005",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3005_ack_0,
          idata => idata,
          odata => tmp821x_xlcssa_3005,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3005
    phi_stmt_3009: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3012_wire;
      req(0) <= phi_stmt_3009_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3009",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3009_ack_0,
          idata => idata,
          odata => conv807x_xlcssa_3009,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3009
    phi_stmt_3140: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3144_wire_constant & type_cast_3146_wire;
      req <= phi_stmt_3140_req_0 & phi_stmt_3140_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3140",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3140_ack_0,
          idata => idata,
          odata => k840x_x1_3140,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3140
    phi_stmt_3147: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3150_wire & type_cast_3152_wire;
      req <= phi_stmt_3147_req_0 & phi_stmt_3147_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3147",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3147_ack_0,
          idata => idata,
          odata => i844x_x2_3147,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3147
    phi_stmt_3153: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3156_wire & type_cast_3159_wire_constant;
      req <= phi_stmt_3153_req_0 & phi_stmt_3153_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3153",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3153_ack_0,
          idata => idata,
          odata => j894x_x1_3153,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3153
    phi_stmt_3558: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3561_wire & type_cast_3564_wire_constant;
      req <= phi_stmt_3558_req_0 & phi_stmt_3558_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3558",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3558_ack_0,
          idata => idata,
          odata => k840x_x0x_xph_3558,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3558
    phi_stmt_3565: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3568_wire & type_cast_3570_wire;
      req <= phi_stmt_3565_req_0 & phi_stmt_3565_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3565",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3565_ack_0,
          idata => idata,
          odata => i844x_x1x_xph_3565,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3565
    phi_stmt_3571: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3574_wire & type_cast_3576_wire;
      req <= phi_stmt_3571_req_0 & phi_stmt_3571_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3571",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3571_ack_0,
          idata => idata,
          odata => j894x_x0x_xph_3571,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3571
    phi_stmt_3580: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3583_wire;
      req(0) <= phi_stmt_3580_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3580",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3580_ack_0,
          idata => idata,
          odata => tmp1040x_xlcssa_3580,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3580
    phi_stmt_3584: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3587_wire;
      req(0) <= phi_stmt_3584_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3584",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3584_ack_0,
          idata => idata,
          odata => conv1025x_xlcssa_3584,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3584
    phi_stmt_3588: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3591_wire;
      req(0) <= phi_stmt_3588_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3588",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3588_ack_0,
          idata => idata,
          odata => tmp1024x_xlcssa_3588,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3588
    phi_stmt_3729: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3732_wire & type_cast_3735_wire_constant;
      req <= phi_stmt_3729_req_0 & phi_stmt_3729_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3729",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3729_ack_0,
          idata => idata,
          odata => k1060x_x1_3729,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3729
    phi_stmt_3736: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3739_wire & type_cast_3741_wire;
      req <= phi_stmt_3736_req_0 & phi_stmt_3736_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3736",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3736_ack_0,
          idata => idata,
          odata => i1068x_x2_3736,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3736
    phi_stmt_3742: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3745_wire & type_cast_3747_wire;
      req <= phi_stmt_3742_req_0 & phi_stmt_3742_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3742",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3742_ack_0,
          idata => idata,
          odata => j1118x_x1_3742,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3742
    phi_stmt_4133: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4136_wire & type_cast_4139_wire_constant;
      req <= phi_stmt_4133_req_0 & phi_stmt_4133_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4133",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4133_ack_0,
          idata => idata,
          odata => k1060x_x0x_xph_4133,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4133
    phi_stmt_4140: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4143_wire & type_cast_4145_wire;
      req <= phi_stmt_4140_req_0 & phi_stmt_4140_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4140",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4140_ack_0,
          idata => idata,
          odata => i1068x_x1x_xph_4140,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4140
    phi_stmt_4146: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4149_wire & type_cast_4151_wire;
      req <= phi_stmt_4146_req_0 & phi_stmt_4146_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4146",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4146_ack_0,
          idata => idata,
          odata => j1118x_x0x_xph_4146,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4146
    phi_stmt_4155: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_4158_wire;
      req(0) <= phi_stmt_4155_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4155",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4155_ack_0,
          idata => idata,
          odata => tmp1262x_xlcssa_4155,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4155
    phi_stmt_4159: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_4162_wire;
      req(0) <= phi_stmt_4159_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4159",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4159_ack_0,
          idata => idata,
          odata => conv1248x_xlcssa_4159,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4159
    phi_stmt_4296: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4300_wire_constant & type_cast_4302_wire;
      req <= phi_stmt_4296_req_0 & phi_stmt_4296_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4296",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4296_ack_0,
          idata => idata,
          odata => k1282x_x1_4296,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4296
    phi_stmt_4303: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4306_wire & type_cast_4308_wire;
      req <= phi_stmt_4303_req_0 & phi_stmt_4303_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4303",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4303_ack_0,
          idata => idata,
          odata => i1286x_x2_4303,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4303
    phi_stmt_4309: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4313_wire_constant & type_cast_4315_wire;
      req <= phi_stmt_4309_req_0 & phi_stmt_4309_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4309",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4309_ack_0,
          idata => idata,
          odata => j1337x_x1_4309,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4309
    phi_stmt_4690: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4694_wire_constant & type_cast_4696_wire;
      req <= phi_stmt_4690_req_0 & phi_stmt_4690_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4690",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4690_ack_0,
          idata => idata,
          odata => k1282x_x0x_xph_4690,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4690
    phi_stmt_4697: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4700_wire & type_cast_4702_wire;
      req <= phi_stmt_4697_req_0 & phi_stmt_4697_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4697",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4697_ack_0,
          idata => idata,
          odata => i1286x_x1x_xph_4697,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4697
    phi_stmt_4703: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4706_wire & type_cast_4708_wire;
      req <= phi_stmt_4703_req_0 & phi_stmt_4703_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4703",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4703_ack_0,
          idata => idata,
          odata => j1337x_x0x_xph_4703,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4703
    phi_stmt_4712: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_4715_wire;
      req(0) <= phi_stmt_4712_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4712",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4712_ack_0,
          idata => idata,
          odata => tmp1481x_xlcssa_4712,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4712
    phi_stmt_4716: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_4719_wire;
      req(0) <= phi_stmt_4716_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4716",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4716_ack_0,
          idata => idata,
          odata => conv1466x_xlcssa_4716,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4716
    phi_stmt_4720: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_4723_wire;
      req(0) <= phi_stmt_4720_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4720",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4720_ack_0,
          idata => idata,
          odata => tmp1465x_xlcssa_4720,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4720
    phi_stmt_4867: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4871_wire_constant & type_cast_4873_wire;
      req <= phi_stmt_4867_req_0 & phi_stmt_4867_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4867",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4867_ack_0,
          idata => idata,
          odata => k1499x_x1_4867,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4867
    phi_stmt_4874: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4877_wire & type_cast_4879_wire;
      req <= phi_stmt_4874_req_0 & phi_stmt_4874_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4874",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4874_ack_0,
          idata => idata,
          odata => i1507x_x2_4874,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4874
    phi_stmt_4880: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4883_wire & type_cast_4885_wire;
      req <= phi_stmt_4880_req_0 & phi_stmt_4880_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4880",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4880_ack_0,
          idata => idata,
          odata => j1558x_x1_4880,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4880
    phi_stmt_5247: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_5250_wire & type_cast_5253_wire_constant;
      req <= phi_stmt_5247_req_0 & phi_stmt_5247_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_5247",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_5247_ack_0,
          idata => idata,
          odata => k1499x_x0x_xph_5247,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_5247
    phi_stmt_5254: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_5257_wire & type_cast_5259_wire;
      req <= phi_stmt_5254_req_0 & phi_stmt_5254_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_5254",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_5254_ack_0,
          idata => idata,
          odata => i1507x_x1x_xph_5254,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_5254
    phi_stmt_5260: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_5263_wire & type_cast_5265_wire;
      req <= phi_stmt_5260_req_0 & phi_stmt_5260_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_5260",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_5260_ack_0,
          idata => idata,
          odata => j1558x_x0x_xph_5260,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_5260
    phi_stmt_899: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_903_wire_constant & type_cast_905_wire;
      req <= phi_stmt_899_req_0 & phi_stmt_899_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_899",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_899_ack_0,
          idata => idata,
          odata => jx_x1_899,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_899
    phi_stmt_906: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_910_wire_constant & type_cast_912_wire;
      req <= phi_stmt_906_req_0 & phi_stmt_906_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_906",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_906_ack_0,
          idata => idata,
          odata => ix_x2_906,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_906
    phi_stmt_913: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_917_wire_constant & type_cast_919_wire;
      req <= phi_stmt_913_req_0 & phi_stmt_913_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_913",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_913_ack_0,
          idata => idata,
          odata => kx_x1_913,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_913
    -- flow-through select operator MUX_1270_inst
    jx_x2_1271 <= type_cast_1268_wire_constant when (cmp160_1255(0) /=  '0') else inc_1227;
    -- flow-through select operator MUX_1820_inst
    j240x_x2_1821 <= div191_1347 when (cmp374_1806(0) /=  '0') else inc365_1784;
    -- flow-through select operator MUX_2383_inst
    j456x_x2_2384 <= type_cast_2381_wire_constant when (cmp592_2368(0) /=  '0') else inc582_2340;
    -- flow-through select operator MUX_2946_inst
    j678x_x2_2947 <= div625_2464 when (cmp812_2932(0) /=  '0') else inc803_2910;
    -- flow-through select operator MUX_3515_inst
    j894x_x2_3516 <= type_cast_3513_wire_constant when (cmp1031_3500(0) /=  '0') else inc1021_3472;
    -- flow-through select operator MUX_4090_inst
    j1118x_x2_4091 <= div1065_3602 when (cmp1253_4076(0) /=  '0') else inc1244_4054;
    -- flow-through select operator MUX_4659_inst
    j1337x_x2_4660 <= type_cast_4657_wire_constant when (cmp1472_4644(0) /=  '0') else inc1462_4616;
    -- flow-through select operator MUX_5216_inst
    j1558x_x2_5217 <= div1504_4734 when (cmp1691_5202(0) /=  '0') else inc1682_5180;
    addr_of_1073_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1073_final_reg_req_0;
      addr_of_1073_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1073_final_reg_req_1;
      addr_of_1073_final_reg_ack_1<= rack(0);
      addr_of_1073_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1073_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1072_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1074,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1156_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1156_final_reg_req_0;
      addr_of_1156_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1156_final_reg_req_1;
      addr_of_1156_final_reg_ack_1<= rack(0);
      addr_of_1156_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1156_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1155_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx131_1157,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1181_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1181_final_reg_req_0;
      addr_of_1181_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1181_final_reg_req_1;
      addr_of_1181_final_reg_ack_1<= rack(0);
      addr_of_1181_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1181_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1180_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx136_1182,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1630_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1630_final_reg_req_0;
      addr_of_1630_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1630_final_reg_req_1;
      addr_of_1630_final_reg_ack_1<= rack(0);
      addr_of_1630_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1630_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1629_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx299_1631,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1713_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1713_final_reg_req_0;
      addr_of_1713_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1713_final_reg_req_1;
      addr_of_1713_final_reg_ack_1<= rack(0);
      addr_of_1713_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1713_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1712_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx342_1714,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1738_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1738_final_reg_req_0;
      addr_of_1738_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1738_final_reg_req_1;
      addr_of_1738_final_reg_ack_1<= rack(0);
      addr_of_1738_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1738_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1737_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx347_1739,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2186_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2186_final_reg_req_0;
      addr_of_2186_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2186_final_reg_req_1;
      addr_of_2186_final_reg_ack_1<= rack(0);
      addr_of_2186_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2186_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2185_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx516_2187,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2269_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2269_final_reg_req_0;
      addr_of_2269_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2269_final_reg_req_1;
      addr_of_2269_final_reg_ack_1<= rack(0);
      addr_of_2269_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2269_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2268_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx559_2270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2294_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2294_final_reg_req_0;
      addr_of_2294_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2294_final_reg_req_1;
      addr_of_2294_final_reg_ack_1<= rack(0);
      addr_of_2294_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2294_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2293_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx564_2295,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2756_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2756_final_reg_req_0;
      addr_of_2756_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2756_final_reg_req_1;
      addr_of_2756_final_reg_ack_1<= rack(0);
      addr_of_2756_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2756_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2755_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx737_2757,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2839_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2839_final_reg_req_0;
      addr_of_2839_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2839_final_reg_req_1;
      addr_of_2839_final_reg_ack_1<= rack(0);
      addr_of_2839_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2839_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2838_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx780_2840,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2864_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2864_final_reg_req_0;
      addr_of_2864_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2864_final_reg_req_1;
      addr_of_2864_final_reg_ack_1<= rack(0);
      addr_of_2864_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2864_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2863_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx785_2865,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3318_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3318_final_reg_req_0;
      addr_of_3318_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3318_final_reg_req_1;
      addr_of_3318_final_reg_ack_1<= rack(0);
      addr_of_3318_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3318_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3317_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx955_3319,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3401_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3401_final_reg_req_0;
      addr_of_3401_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3401_final_reg_req_1;
      addr_of_3401_final_reg_ack_1<= rack(0);
      addr_of_3401_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3401_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3400_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx998_3402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3426_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3426_final_reg_req_0;
      addr_of_3426_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3426_final_reg_req_1;
      addr_of_3426_final_reg_ack_1<= rack(0);
      addr_of_3426_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3426_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3425_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1003_3427,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3900_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3900_final_reg_req_0;
      addr_of_3900_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3900_final_reg_req_1;
      addr_of_3900_final_reg_ack_1<= rack(0);
      addr_of_3900_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3900_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3899_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1178_3901,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3983_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3983_final_reg_req_0;
      addr_of_3983_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3983_final_reg_req_1;
      addr_of_3983_final_reg_ack_1<= rack(0);
      addr_of_3983_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3983_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3982_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1221_3984,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4008_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4008_final_reg_req_0;
      addr_of_4008_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4008_final_reg_req_1;
      addr_of_4008_final_reg_ack_1<= rack(0);
      addr_of_4008_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4008_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4007_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1226_4009,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4462_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4462_final_reg_req_0;
      addr_of_4462_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4462_final_reg_req_1;
      addr_of_4462_final_reg_ack_1<= rack(0);
      addr_of_4462_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4462_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4461_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1396_4463,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4545_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4545_final_reg_req_0;
      addr_of_4545_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4545_final_reg_req_1;
      addr_of_4545_final_reg_ack_1<= rack(0);
      addr_of_4545_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4545_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4544_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1439_4546,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4570_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4570_final_reg_req_0;
      addr_of_4570_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4570_final_reg_req_1;
      addr_of_4570_final_reg_ack_1<= rack(0);
      addr_of_4570_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4570_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4569_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1444_4571,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_5026_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_5026_final_reg_req_0;
      addr_of_5026_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_5026_final_reg_req_1;
      addr_of_5026_final_reg_ack_1<= rack(0);
      addr_of_5026_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_5026_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_5025_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1616_5027,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_5109_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_5109_final_reg_req_0;
      addr_of_5109_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_5109_final_reg_req_1;
      addr_of_5109_final_reg_ack_1<= rack(0);
      addr_of_5109_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_5109_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_5108_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1659_5110,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_5134_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_5134_final_reg_req_0;
      addr_of_5134_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_5134_final_reg_req_1;
      addr_of_5134_final_reg_ack_1<= rack(0);
      addr_of_5134_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_5134_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_5133_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1664_5135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1011_inst
    process(conv60_976) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv60_976(31 downto 0);
      type_cast_1011_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1013_inst
    process(add73_1008) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add73_1008(31 downto 0);
      type_cast_1013_wire <= tmp_var; -- 
    end process;
    type_cast_1026_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1026_inst_req_0;
      type_cast_1026_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1026_inst_req_1;
      type_cast_1026_inst_ack_1<= rack(0);
      type_cast_1026_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1026_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1025_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_1027,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1031_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1031_inst_req_0;
      type_cast_1031_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1031_inst_req_1;
      type_cast_1031_inst_ack_1<= rack(0);
      type_cast_1031_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1031_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1030_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_1032,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1055_inst
    process(add90_1052) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add90_1052(31 downto 0);
      type_cast_1055_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1060_inst
    process(ASHR_i32_i32_1059_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1059_wire(31 downto 0);
      shr_1061 <= tmp_var; -- 
    end process;
    type_cast_1066_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1066_inst_req_0;
      type_cast_1066_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1066_inst_req_1;
      type_cast_1066_inst_ack_1<= rack(0);
      type_cast_1066_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1066_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1065_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1067,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1085_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1085_inst_req_0;
      type_cast_1085_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1085_inst_req_1;
      type_cast_1085_inst_ack_1<= rack(0);
      type_cast_1085_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1085_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1084_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1086,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1139_inst
    process(add111_1116) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add111_1116(31 downto 0);
      type_cast_1139_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1144_inst
    process(ASHR_i32_i32_1143_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1143_wire(31 downto 0);
      shr129_1145 <= tmp_var; -- 
    end process;
    type_cast_1149_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1149_inst_req_0;
      type_cast_1149_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1149_inst_req_1;
      type_cast_1149_inst_ack_1<= rack(0);
      type_cast_1149_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1149_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1148_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom130_1150,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1164_inst
    process(add127_1136) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add127_1136(31 downto 0);
      type_cast_1164_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1169_inst
    process(ASHR_i32_i32_1168_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1168_wire(31 downto 0);
      shr134_1170 <= tmp_var; -- 
    end process;
    type_cast_1174_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1174_inst_req_0;
      type_cast_1174_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1174_inst_req_1;
      type_cast_1174_inst_ack_1<= rack(0);
      type_cast_1174_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1174_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1173_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom135_1175,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1192_inst_req_0;
      type_cast_1192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1192_inst_req_1;
      type_cast_1192_inst_ack_1<= rack(0);
      type_cast_1192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1191_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv139_1193,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1202_inst
    process(add140_1199) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add140_1199(31 downto 0);
      type_cast_1202_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1204_inst
    process(conv31_811) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv31_811(31 downto 0);
      type_cast_1204_wire <= tmp_var; -- 
    end process;
    type_cast_1231_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1231_inst_req_0;
      type_cast_1231_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1231_inst_req_1;
      type_cast_1231_inst_ack_1<= rack(0);
      type_cast_1231_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1231_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1230_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_1232,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp154_1235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1258_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1258_inst_req_0;
      type_cast_1258_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1258_inst_req_1;
      type_cast_1258_inst_ack_1<= rack(0);
      type_cast_1258_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1258_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp160_1255,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc165_1259,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1275_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1275_inst_req_0;
      type_cast_1275_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1275_inst_req_1;
      type_cast_1275_inst_ack_1<= rack(0);
      type_cast_1275_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1275_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1274_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv168_1276,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1282_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1282_inst_req_0;
      type_cast_1282_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1282_inst_req_1;
      type_cast_1282_inst_ack_1<= rack(0);
      type_cast_1282_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1282_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp169_1279,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1283,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1310_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1310_inst_req_0;
      type_cast_1310_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1310_inst_req_1;
      type_cast_1310_inst_ack_1<= rack(0);
      type_cast_1310_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1310_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_1271,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1310_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1312_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1312_inst_req_0;
      type_cast_1312_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1312_inst_req_1;
      type_cast_1312_inst_ack_1<= rack(0);
      type_cast_1312_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1312_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_899,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1312_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1316_inst_req_0;
      type_cast_1316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1316_inst_req_1;
      type_cast_1316_inst_ack_1<= rack(0);
      type_cast_1316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1316_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_906,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1316_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1318_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1318_inst_req_0;
      type_cast_1318_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1318_inst_req_1;
      type_cast_1318_inst_ack_1<= rack(0);
      type_cast_1318_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1318_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc165x_xix_x2_1264,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1318_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1325_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1325_inst_req_0;
      type_cast_1325_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1325_inst_req_1;
      type_cast_1325_inst_ack_1<= rack(0);
      type_cast_1325_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1325_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add148_1219,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1325_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1332_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1332_inst_req_0;
      type_cast_1332_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1332_inst_req_1;
      type_cast_1332_inst_ack_1<= rack(0);
      type_cast_1332_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1332_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv155_1239,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1332_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1336_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1336_inst_req_0;
      type_cast_1336_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1336_inst_req_1;
      type_cast_1336_inst_ack_1<= rack(0);
      type_cast_1336_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1336_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp154_1235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1336_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1340_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1340_inst_req_0;
      type_cast_1340_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1340_inst_req_1;
      type_cast_1340_inst_ack_1<= rack(0);
      type_cast_1340_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1340_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp154x_xlcssa_1333,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv190_1341,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1380_inst_req_0;
      type_cast_1380_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1380_inst_req_1;
      type_cast_1380_inst_ack_1<= rack(0);
      type_cast_1380_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1380_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp201_1353,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv226_1381,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1390_inst
    process(sext1766_1387) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1766_1387(31 downto 0);
      type_cast_1390_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1395_inst
    process(ASHR_i32_i32_1394_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1394_wire(31 downto 0);
      conv234_1396 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1405_inst
    process(sext1718_1402) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1718_1402(31 downto 0);
      type_cast_1405_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1410_inst
    process(ASHR_i32_i32_1409_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1409_wire(31 downto 0);
      conv236_1411 <= tmp_var; -- 
    end process;
    type_cast_1419_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1419_inst_req_0;
      type_cast_1419_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1419_inst_req_1;
      type_cast_1419_inst_ack_1<= rack(0);
      type_cast_1419_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1419_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp197_1350,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv248_1420,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1429_inst
    process(sext1767_1426) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1767_1426(31 downto 0);
      type_cast_1429_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1434_inst
    process(ASHR_i32_i32_1433_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1433_wire(31 downto 0);
      conv291_1435 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1455_inst
    process(sext1719_1452) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1719_1452(31 downto 0);
      type_cast_1455_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1460_inst
    process(ASHR_i32_i32_1459_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1459_wire(31 downto 0);
      conv315_1461 <= tmp_var; -- 
    end process;
    type_cast_1467_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1467_inst_req_0;
      type_cast_1467_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1467_inst_req_1;
      type_cast_1467_inst_ack_1<= rack(0);
      type_cast_1467_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1467_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div191_1347,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1467_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1469_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1469_inst_req_0;
      type_cast_1469_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1469_inst_req_1;
      type_cast_1469_inst_ack_1<= rack(0);
      type_cast_1469_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1469_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j240x_x0x_xph_1857,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1469_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1476_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1476_inst_req_0;
      type_cast_1476_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1476_inst_req_1;
      type_cast_1476_inst_ack_1<= rack(0);
      type_cast_1476_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1476_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i194x_x1x_xph_1863,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1476_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1483_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1483_inst_req_0;
      type_cast_1483_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1483_inst_req_1;
      type_cast_1483_inst_ack_1<= rack(0);
      type_cast_1483_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1483_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k186x_x0x_xph_1869,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1483_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1488_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1488_inst_req_0;
      type_cast_1488_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1488_inst_req_1;
      type_cast_1488_inst_ack_1<= rack(0);
      type_cast_1488_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1488_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1487_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv246_1489,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1492_inst
    process(conv246_1489) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv246_1489(31 downto 0);
      type_cast_1492_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1494_inst
    process(conv248_1420) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv248_1420(31 downto 0);
      type_cast_1494_wire <= tmp_var; -- 
    end process;
    type_cast_1509_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1509_inst_req_0;
      type_cast_1509_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1509_inst_req_1;
      type_cast_1509_inst_ack_1<= rack(0);
      type_cast_1509_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1509_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp254_1506,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_1510,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1524_inst
    process(conv246_1489) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv246_1489(31 downto 0);
      type_cast_1524_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1526_inst
    process(add259_1521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add259_1521(31 downto 0);
      type_cast_1526_wire <= tmp_var; -- 
    end process;
    type_cast_1539_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1539_inst_req_0;
      type_cast_1539_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1539_inst_req_1;
      type_cast_1539_inst_ack_1<= rack(0);
      type_cast_1539_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1539_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1538_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv264_1540,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1543_inst
    process(conv264_1540) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv264_1540(31 downto 0);
      type_cast_1543_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1545_inst
    process(conv248_1420) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv248_1420(31 downto 0);
      type_cast_1545_wire <= tmp_var; -- 
    end process;
    type_cast_1560_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1560_inst_req_0;
      type_cast_1560_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1560_inst_req_1;
      type_cast_1560_inst_ack_1<= rack(0);
      type_cast_1560_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1560_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp272_1557,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv273_1561,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1569_inst
    process(conv264_1540) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv264_1540(31 downto 0);
      type_cast_1569_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1571_inst
    process(add276_1566) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add276_1566(31 downto 0);
      type_cast_1571_wire <= tmp_var; -- 
    end process;
    type_cast_1584_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1584_inst_req_0;
      type_cast_1584_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1584_inst_req_1;
      type_cast_1584_inst_ack_1<= rack(0);
      type_cast_1584_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1584_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1583_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv283_1585,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1589_inst_req_0;
      type_cast_1589_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1589_inst_req_1;
      type_cast_1589_inst_ack_1<= rack(0);
      type_cast_1589_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1589_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1588_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv287_1590,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1613_inst
    process(add295_1610) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add295_1610(31 downto 0);
      type_cast_1613_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1618_inst
    process(ASHR_i32_i32_1617_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1617_wire(31 downto 0);
      shr297_1619 <= tmp_var; -- 
    end process;
    type_cast_1623_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1623_inst_req_0;
      type_cast_1623_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1623_inst_req_1;
      type_cast_1623_inst_ack_1<= rack(0);
      type_cast_1623_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1623_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1622_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom298_1624,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1642_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1642_inst_req_0;
      type_cast_1642_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1642_inst_req_1;
      type_cast_1642_inst_ack_1<= rack(0);
      type_cast_1642_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1642_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1641_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv304_1643,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1696_inst
    process(add322_1673) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add322_1673(31 downto 0);
      type_cast_1696_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1701_inst
    process(ASHR_i32_i32_1700_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1700_wire(31 downto 0);
      shr340_1702 <= tmp_var; -- 
    end process;
    type_cast_1706_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1706_inst_req_0;
      type_cast_1706_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1706_inst_req_1;
      type_cast_1706_inst_ack_1<= rack(0);
      type_cast_1706_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1706_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1705_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom341_1707,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1721_inst
    process(add338_1693) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add338_1693(31 downto 0);
      type_cast_1721_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1726_inst
    process(ASHR_i32_i32_1725_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1725_wire(31 downto 0);
      shr345_1727 <= tmp_var; -- 
    end process;
    type_cast_1731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1731_inst_req_0;
      type_cast_1731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1731_inst_req_1;
      type_cast_1731_inst_ack_1<= rack(0);
      type_cast_1731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1731_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1730_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom346_1732,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1749_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1749_inst_req_0;
      type_cast_1749_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1749_inst_req_1;
      type_cast_1749_inst_ack_1<= rack(0);
      type_cast_1749_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1749_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1748_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv352_1750,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1759_inst
    process(add353_1756) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add353_1756(31 downto 0);
      type_cast_1759_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1761_inst
    process(conv226_1381) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv226_1381(31 downto 0);
      type_cast_1761_wire <= tmp_var; -- 
    end process;
    type_cast_1788_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1788_inst_req_0;
      type_cast_1788_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1788_inst_req_1;
      type_cast_1788_inst_ack_1<= rack(0);
      type_cast_1788_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1788_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1787_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv367_1789,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1795_inst_req_0;
      type_cast_1795_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1795_inst_req_1;
      type_cast_1795_inst_ack_1<= rack(0);
      type_cast_1795_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1795_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp368_1792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv369_1796,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1809_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1809_inst_req_0;
      type_cast_1809_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1809_inst_req_1;
      type_cast_1809_inst_ack_1<= rack(0);
      type_cast_1809_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1809_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp374_1806,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc379_1810,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1825_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1825_inst_req_0;
      type_cast_1825_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1825_inst_req_1;
      type_cast_1825_inst_ack_1<= rack(0);
      type_cast_1825_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1825_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1824_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv382_1826,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1832_inst_req_0;
      type_cast_1832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1832_inst_req_1;
      type_cast_1832_inst_ack_1<= rack(0);
      type_cast_1832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1832_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp383_1829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv384_1833,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1860_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1860_inst_req_0;
      type_cast_1860_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1860_inst_req_1;
      type_cast_1860_inst_ack_1<= rack(0);
      type_cast_1860_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1860_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j240x_x1_1464,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1860_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1862_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1862_inst_req_0;
      type_cast_1862_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1862_inst_req_1;
      type_cast_1862_inst_ack_1<= rack(0);
      type_cast_1862_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1862_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j240x_x2_1821,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1862_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1866_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1866_inst_req_0;
      type_cast_1866_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1866_inst_req_1;
      type_cast_1866_inst_ack_1<= rack(0);
      type_cast_1866_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1866_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i194x_x2_1470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1866_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1868_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1868_inst_req_0;
      type_cast_1868_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1868_inst_req_1;
      type_cast_1868_inst_ack_1<= rack(0);
      type_cast_1868_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1868_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc379x_xi194x_x2_1815,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1868_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1872_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1872_inst_req_0;
      type_cast_1872_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1872_inst_req_1;
      type_cast_1872_inst_ack_1<= rack(0);
      type_cast_1872_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1872_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add361_1776,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1872_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1882_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1882_inst_req_0;
      type_cast_1882_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1882_inst_req_1;
      type_cast_1882_inst_ack_1<= rack(0);
      type_cast_1882_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1882_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp383_1829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1882_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1886_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1886_inst_req_0;
      type_cast_1886_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1886_inst_req_1;
      type_cast_1886_inst_ack_1<= rack(0);
      type_cast_1886_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1886_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv369_1796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1886_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1890_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1890_inst_req_0;
      type_cast_1890_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1890_inst_req_1;
      type_cast_1890_inst_ack_1<= rack(0);
      type_cast_1890_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1890_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp383x_xlcssa_1879,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv408_1891,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1930_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1930_inst_req_0;
      type_cast_1930_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1930_inst_req_1;
      type_cast_1930_inst_ack_1<= rack(0);
      type_cast_1930_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1930_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp417_1903,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv442_1931,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1940_inst
    process(sext1768_1937) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1768_1937(31 downto 0);
      type_cast_1940_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1945_inst
    process(ASHR_i32_i32_1944_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1944_wire(31 downto 0);
      conv450_1946 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1955_inst
    process(sext1720_1952) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1720_1952(31 downto 0);
      type_cast_1955_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1960_inst
    process(ASHR_i32_i32_1959_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1959_wire(31 downto 0);
      conv452_1961 <= tmp_var; -- 
    end process;
    type_cast_1969_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1969_inst_req_0;
      type_cast_1969_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1969_inst_req_1;
      type_cast_1969_inst_ack_1<= rack(0);
      type_cast_1969_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1969_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp413_1900,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv464_1970,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1979_inst
    process(sext1769_1976) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1769_1976(31 downto 0);
      type_cast_1979_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1984_inst
    process(ASHR_i32_i32_1983_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1983_wire(31 downto 0);
      conv508_1985 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2005_inst
    process(sext1721_2002) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1721_2002(31 downto 0);
      type_cast_2005_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2010_inst
    process(ASHR_i32_i32_2009_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2009_wire(31 downto 0);
      conv532_2011 <= tmp_var; -- 
    end process;
    type_cast_2017_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2017_inst_req_0;
      type_cast_2017_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2017_inst_req_1;
      type_cast_2017_inst_ack_1<= rack(0);
      type_cast_2017_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2017_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k402x_x0x_xph_2420,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2017_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2024_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2024_inst_req_0;
      type_cast_2024_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2024_inst_req_1;
      type_cast_2024_inst_ack_1<= rack(0);
      type_cast_2024_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2024_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div409_1897,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2024_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2026_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2026_inst_req_0;
      type_cast_2026_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2026_inst_req_1;
      type_cast_2026_inst_ack_1<= rack(0);
      type_cast_2026_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2026_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i406x_x1x_xph_2427,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2026_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2030_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2030_inst_req_0;
      type_cast_2030_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2030_inst_req_1;
      type_cast_2030_inst_ack_1<= rack(0);
      type_cast_2030_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2030_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j456x_x0x_xph_2433,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2030_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2038_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2038_inst_req_0;
      type_cast_2038_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2038_inst_req_1;
      type_cast_2038_inst_ack_1<= rack(0);
      type_cast_2038_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2038_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2037_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv462_2039,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2042_inst
    process(conv462_2039) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv462_2039(31 downto 0);
      type_cast_2042_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2044_inst
    process(conv464_1970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv464_1970(31 downto 0);
      type_cast_2044_wire <= tmp_var; -- 
    end process;
    type_cast_2059_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2059_inst_req_0;
      type_cast_2059_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2059_inst_req_1;
      type_cast_2059_inst_ack_1<= rack(0);
      type_cast_2059_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2059_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp470_2056,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv471_2060,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2074_inst
    process(conv462_2039) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv462_2039(31 downto 0);
      type_cast_2074_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2076_inst
    process(add475_2071) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add475_2071(31 downto 0);
      type_cast_2076_wire <= tmp_var; -- 
    end process;
    type_cast_2089_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2089_inst_req_0;
      type_cast_2089_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2089_inst_req_1;
      type_cast_2089_inst_ack_1<= rack(0);
      type_cast_2089_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2089_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2088_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv480_2090,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2093_inst
    process(conv480_2090) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv480_2090(31 downto 0);
      type_cast_2093_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2095_inst
    process(conv464_1970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv464_1970(31 downto 0);
      type_cast_2095_wire <= tmp_var; -- 
    end process;
    type_cast_2110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2110_inst_req_0;
      type_cast_2110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2110_inst_req_1;
      type_cast_2110_inst_ack_1<= rack(0);
      type_cast_2110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp488_2107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv489_2111,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2125_inst
    process(conv480_2090) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv480_2090(31 downto 0);
      type_cast_2125_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2127_inst
    process(add493_2122) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add493_2122(31 downto 0);
      type_cast_2127_wire <= tmp_var; -- 
    end process;
    type_cast_2140_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2140_inst_req_0;
      type_cast_2140_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2140_inst_req_1;
      type_cast_2140_inst_ack_1<= rack(0);
      type_cast_2140_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2140_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2139_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv500_2141,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2145_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2145_inst_req_0;
      type_cast_2145_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2145_inst_req_1;
      type_cast_2145_inst_ack_1<= rack(0);
      type_cast_2145_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2145_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2144_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv504_2146,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2169_inst
    process(add512_2166) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add512_2166(31 downto 0);
      type_cast_2169_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2174_inst
    process(ASHR_i32_i32_2173_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2173_wire(31 downto 0);
      shr514_2175 <= tmp_var; -- 
    end process;
    type_cast_2179_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2179_inst_req_0;
      type_cast_2179_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2179_inst_req_1;
      type_cast_2179_inst_ack_1<= rack(0);
      type_cast_2179_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2179_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2178_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom515_2180,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2198_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2198_inst_req_0;
      type_cast_2198_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2198_inst_req_1;
      type_cast_2198_inst_ack_1<= rack(0);
      type_cast_2198_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2198_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2197_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv521_2199,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2252_inst
    process(add539_2229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add539_2229(31 downto 0);
      type_cast_2252_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2257_inst
    process(ASHR_i32_i32_2256_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2256_wire(31 downto 0);
      shr557_2258 <= tmp_var; -- 
    end process;
    type_cast_2262_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2262_inst_req_0;
      type_cast_2262_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2262_inst_req_1;
      type_cast_2262_inst_ack_1<= rack(0);
      type_cast_2262_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2262_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2261_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom558_2263,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2277_inst
    process(add555_2249) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add555_2249(31 downto 0);
      type_cast_2277_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2282_inst
    process(ASHR_i32_i32_2281_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2281_wire(31 downto 0);
      shr562_2283 <= tmp_var; -- 
    end process;
    type_cast_2287_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2287_inst_req_0;
      type_cast_2287_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2287_inst_req_1;
      type_cast_2287_inst_ack_1<= rack(0);
      type_cast_2287_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2287_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2286_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom563_2288,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2305_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2305_inst_req_0;
      type_cast_2305_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2305_inst_req_1;
      type_cast_2305_inst_ack_1<= rack(0);
      type_cast_2305_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2305_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2304_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv569_2306,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2315_inst
    process(add570_2312) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add570_2312(31 downto 0);
      type_cast_2315_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2317_inst
    process(conv442_1931) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv442_1931(31 downto 0);
      type_cast_2317_wire <= tmp_var; -- 
    end process;
    type_cast_2344_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2344_inst_req_0;
      type_cast_2344_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2344_inst_req_1;
      type_cast_2344_inst_ack_1<= rack(0);
      type_cast_2344_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2344_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2343_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv584_2345,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2351_inst_req_0;
      type_cast_2351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2351_inst_req_1;
      type_cast_2351_inst_ack_1<= rack(0);
      type_cast_2351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp585_2348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv586_2352,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2371_inst_req_0;
      type_cast_2371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2371_inst_req_1;
      type_cast_2371_inst_ack_1<= rack(0);
      type_cast_2371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp592_2368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc597_2372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2388_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2388_inst_req_0;
      type_cast_2388_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2388_inst_req_1;
      type_cast_2388_inst_ack_1<= rack(0);
      type_cast_2388_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2388_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2387_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv600_2389,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2395_inst_req_0;
      type_cast_2395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2395_inst_req_1;
      type_cast_2395_inst_ack_1<= rack(0);
      type_cast_2395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp601_2392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv602_2396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2423_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2423_inst_req_0;
      type_cast_2423_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2423_inst_req_1;
      type_cast_2423_inst_ack_1<= rack(0);
      type_cast_2423_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2423_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add578_2332,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2423_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2430_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2430_inst_req_0;
      type_cast_2430_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2430_inst_req_1;
      type_cast_2430_inst_ack_1<= rack(0);
      type_cast_2430_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2430_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i406x_x2_2021,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2430_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2432_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2432_inst_req_0;
      type_cast_2432_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2432_inst_req_1;
      type_cast_2432_inst_ack_1<= rack(0);
      type_cast_2432_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2432_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc597x_xi406x_x2_2377,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2432_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2436_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2436_inst_req_0;
      type_cast_2436_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2436_inst_req_1;
      type_cast_2436_inst_ack_1<= rack(0);
      type_cast_2436_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2436_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j456x_x1_2027,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2436_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2438_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2438_inst_req_0;
      type_cast_2438_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2438_inst_req_1;
      type_cast_2438_inst_ack_1<= rack(0);
      type_cast_2438_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2438_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j456x_x2_2384,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2438_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2445_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2445_inst_req_0;
      type_cast_2445_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2445_inst_req_1;
      type_cast_2445_inst_ack_1<= rack(0);
      type_cast_2445_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2445_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp601_2392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2445_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2449_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2449_inst_req_0;
      type_cast_2449_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2449_inst_req_1;
      type_cast_2449_inst_ack_1<= rack(0);
      type_cast_2449_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2449_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv586_2352,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2449_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2453_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2453_inst_req_0;
      type_cast_2453_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2453_inst_req_1;
      type_cast_2453_inst_ack_1<= rack(0);
      type_cast_2453_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2453_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp585_2348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2453_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2457_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2457_inst_req_0;
      type_cast_2457_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2457_inst_req_1;
      type_cast_2457_inst_ack_1<= rack(0);
      type_cast_2457_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2457_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp585x_xlcssa_2450,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv624_2458,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2467_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2467_inst_req_0;
      type_cast_2467_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2467_inst_req_1;
      type_cast_2467_inst_ack_1<= rack(0);
      type_cast_2467_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2467_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp601x_xlcssa_2442,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv630_2468,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2507_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2507_inst_req_0;
      type_cast_2507_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2507_inst_req_1;
      type_cast_2507_inst_ack_1<= rack(0);
      type_cast_2507_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2507_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp639_2480,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv664_2508,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2517_inst
    process(sext1770_2514) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1770_2514(31 downto 0);
      type_cast_2517_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2522_inst
    process(ASHR_i32_i32_2521_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2521_wire(31 downto 0);
      conv672_2523 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2532_inst
    process(sext1722_2529) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1722_2529(31 downto 0);
      type_cast_2532_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2537_inst
    process(ASHR_i32_i32_2536_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2536_wire(31 downto 0);
      conv674_2538 <= tmp_var; -- 
    end process;
    type_cast_2546_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2546_inst_req_0;
      type_cast_2546_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2546_inst_req_1;
      type_cast_2546_inst_ack_1<= rack(0);
      type_cast_2546_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2546_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp635_2477,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv686_2547,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2556_inst
    process(sext1771_2553) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1771_2553(31 downto 0);
      type_cast_2556_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2561_inst
    process(ASHR_i32_i32_2560_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2560_wire(31 downto 0);
      conv729_2562 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2582_inst
    process(sext1723_2579) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1723_2579(31 downto 0);
      type_cast_2582_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2587_inst
    process(ASHR_i32_i32_2586_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2586_wire(31 downto 0);
      conv753_2588 <= tmp_var; -- 
    end process;
    type_cast_2597_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2597_inst_req_0;
      type_cast_2597_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2597_inst_req_1;
      type_cast_2597_inst_ack_1<= rack(0);
      type_cast_2597_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2597_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k620x_x0x_xph_2983,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2597_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2601_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2601_inst_req_0;
      type_cast_2601_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2601_inst_req_1;
      type_cast_2601_inst_ack_1<= rack(0);
      type_cast_2601_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2601_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div631_2474,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2601_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2603_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2603_inst_req_0;
      type_cast_2603_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2603_inst_req_1;
      type_cast_2603_inst_ack_1<= rack(0);
      type_cast_2603_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2603_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i628x_x1x_xph_2990,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2603_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2607_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2607_inst_req_0;
      type_cast_2607_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2607_inst_req_1;
      type_cast_2607_inst_ack_1<= rack(0);
      type_cast_2607_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2607_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div625_2464,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2607_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2609_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2609_inst_req_0;
      type_cast_2609_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2609_inst_req_1;
      type_cast_2609_inst_ack_1<= rack(0);
      type_cast_2609_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2609_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j678x_x0x_xph_2996,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2609_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2614_inst_req_0;
      type_cast_2614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2614_inst_req_1;
      type_cast_2614_inst_ack_1<= rack(0);
      type_cast_2614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2613_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv684_2615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2618_inst
    process(conv684_2615) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv684_2615(31 downto 0);
      type_cast_2618_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2620_inst
    process(conv686_2547) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv686_2547(31 downto 0);
      type_cast_2620_wire <= tmp_var; -- 
    end process;
    type_cast_2635_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2635_inst_req_0;
      type_cast_2635_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2635_inst_req_1;
      type_cast_2635_inst_ack_1<= rack(0);
      type_cast_2635_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2635_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp692_2632,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv693_2636,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2650_inst
    process(conv684_2615) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv684_2615(31 downto 0);
      type_cast_2650_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2652_inst
    process(add697_2647) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add697_2647(31 downto 0);
      type_cast_2652_wire <= tmp_var; -- 
    end process;
    type_cast_2665_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2665_inst_req_0;
      type_cast_2665_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2665_inst_req_1;
      type_cast_2665_inst_ack_1<= rack(0);
      type_cast_2665_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2665_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2664_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv702_2666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2669_inst
    process(conv702_2666) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv702_2666(31 downto 0);
      type_cast_2669_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2671_inst
    process(conv686_2547) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv686_2547(31 downto 0);
      type_cast_2671_wire <= tmp_var; -- 
    end process;
    type_cast_2686_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2686_inst_req_0;
      type_cast_2686_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2686_inst_req_1;
      type_cast_2686_inst_ack_1<= rack(0);
      type_cast_2686_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2686_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp710_2683,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv711_2687,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2695_inst
    process(conv702_2666) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv702_2666(31 downto 0);
      type_cast_2695_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2697_inst
    process(add714_2692) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add714_2692(31 downto 0);
      type_cast_2697_wire <= tmp_var; -- 
    end process;
    type_cast_2710_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2710_inst_req_0;
      type_cast_2710_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2710_inst_req_1;
      type_cast_2710_inst_ack_1<= rack(0);
      type_cast_2710_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2710_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2709_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv721_2711,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2715_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2715_inst_req_0;
      type_cast_2715_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2715_inst_req_1;
      type_cast_2715_inst_ack_1<= rack(0);
      type_cast_2715_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2715_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2714_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv725_2716,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2739_inst
    process(add733_2736) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add733_2736(31 downto 0);
      type_cast_2739_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2744_inst
    process(ASHR_i32_i32_2743_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2743_wire(31 downto 0);
      shr735_2745 <= tmp_var; -- 
    end process;
    type_cast_2749_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2749_inst_req_0;
      type_cast_2749_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2749_inst_req_1;
      type_cast_2749_inst_ack_1<= rack(0);
      type_cast_2749_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2749_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2748_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom736_2750,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2768_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2768_inst_req_0;
      type_cast_2768_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2768_inst_req_1;
      type_cast_2768_inst_ack_1<= rack(0);
      type_cast_2768_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2768_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2767_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv742_2769,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2822_inst
    process(add760_2799) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add760_2799(31 downto 0);
      type_cast_2822_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2827_inst
    process(ASHR_i32_i32_2826_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2826_wire(31 downto 0);
      shr778_2828 <= tmp_var; -- 
    end process;
    type_cast_2832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2832_inst_req_0;
      type_cast_2832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2832_inst_req_1;
      type_cast_2832_inst_ack_1<= rack(0);
      type_cast_2832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2832_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2831_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom779_2833,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2847_inst
    process(add776_2819) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add776_2819(31 downto 0);
      type_cast_2847_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2852_inst
    process(ASHR_i32_i32_2851_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2851_wire(31 downto 0);
      shr783_2853 <= tmp_var; -- 
    end process;
    type_cast_2857_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2857_inst_req_0;
      type_cast_2857_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2857_inst_req_1;
      type_cast_2857_inst_ack_1<= rack(0);
      type_cast_2857_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2857_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2856_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom784_2858,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2875_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2875_inst_req_0;
      type_cast_2875_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2875_inst_req_1;
      type_cast_2875_inst_ack_1<= rack(0);
      type_cast_2875_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2875_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2874_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv790_2876,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2885_inst
    process(add791_2882) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add791_2882(31 downto 0);
      type_cast_2885_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2887_inst
    process(conv664_2508) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv664_2508(31 downto 0);
      type_cast_2887_wire <= tmp_var; -- 
    end process;
    type_cast_2914_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2914_inst_req_0;
      type_cast_2914_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2914_inst_req_1;
      type_cast_2914_inst_ack_1<= rack(0);
      type_cast_2914_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2914_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2913_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv805_2915,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2921_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2921_inst_req_0;
      type_cast_2921_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2921_inst_req_1;
      type_cast_2921_inst_ack_1<= rack(0);
      type_cast_2921_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2921_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp806_2918,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv807_2922,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2935_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2935_inst_req_0;
      type_cast_2935_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2935_inst_req_1;
      type_cast_2935_inst_ack_1<= rack(0);
      type_cast_2935_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2935_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp812_2932,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc817_2936,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2951_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2951_inst_req_0;
      type_cast_2951_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2951_inst_req_1;
      type_cast_2951_inst_ack_1<= rack(0);
      type_cast_2951_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2951_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2950_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv820_2952,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2958_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2958_inst_req_0;
      type_cast_2958_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2958_inst_req_1;
      type_cast_2958_inst_ack_1<= rack(0);
      type_cast_2958_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2958_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp821_2955,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv822_2959,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2986_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2986_inst_req_0;
      type_cast_2986_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2986_inst_req_1;
      type_cast_2986_inst_ack_1<= rack(0);
      type_cast_2986_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2986_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add799_2902,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2986_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2993_inst_req_0;
      type_cast_2993_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2993_inst_req_1;
      type_cast_2993_inst_ack_1<= rack(0);
      type_cast_2993_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2993_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i628x_x2_2598,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2993_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2995_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2995_inst_req_0;
      type_cast_2995_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2995_inst_req_1;
      type_cast_2995_inst_ack_1<= rack(0);
      type_cast_2995_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2995_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc817x_xi628x_x2_2941,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2995_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2999_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2999_inst_req_0;
      type_cast_2999_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2999_inst_req_1;
      type_cast_2999_inst_ack_1<= rack(0);
      type_cast_2999_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2999_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j678x_x1_2604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2999_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3001_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3001_inst_req_0;
      type_cast_3001_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3001_inst_req_1;
      type_cast_3001_inst_ack_1<= rack(0);
      type_cast_3001_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3001_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j678x_x2_2947,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3001_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3008_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3008_inst_req_0;
      type_cast_3008_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3008_inst_req_1;
      type_cast_3008_inst_ack_1<= rack(0);
      type_cast_3008_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3008_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp821_2955,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3008_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3012_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3012_inst_req_0;
      type_cast_3012_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3012_inst_req_1;
      type_cast_3012_inst_ack_1<= rack(0);
      type_cast_3012_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3012_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv807_2922,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3012_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3016_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3016_inst_req_0;
      type_cast_3016_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3016_inst_req_1;
      type_cast_3016_inst_ack_1<= rack(0);
      type_cast_3016_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3016_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp821x_xlcssa_3005,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv846_3017,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3056_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3056_inst_req_0;
      type_cast_3056_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3056_inst_req_1;
      type_cast_3056_inst_ack_1<= rack(0);
      type_cast_3056_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3056_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp855_3029,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv880_3057,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3066_inst
    process(sext1772_3063) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1772_3063(31 downto 0);
      type_cast_3066_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3071_inst
    process(ASHR_i32_i32_3070_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3070_wire(31 downto 0);
      conv888_3072 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3081_inst
    process(sext1724_3078) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1724_3078(31 downto 0);
      type_cast_3081_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3086_inst
    process(ASHR_i32_i32_3085_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3085_wire(31 downto 0);
      conv890_3087 <= tmp_var; -- 
    end process;
    type_cast_3095_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3095_inst_req_0;
      type_cast_3095_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3095_inst_req_1;
      type_cast_3095_inst_ack_1<= rack(0);
      type_cast_3095_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3095_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp851_3026,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv902_3096,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3105_inst
    process(sext1773_3102) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1773_3102(31 downto 0);
      type_cast_3105_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3110_inst
    process(ASHR_i32_i32_3109_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3109_wire(31 downto 0);
      conv947_3111 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3131_inst
    process(sext1725_3128) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1725_3128(31 downto 0);
      type_cast_3131_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3136_inst
    process(ASHR_i32_i32_3135_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3135_wire(31 downto 0);
      conv971_3137 <= tmp_var; -- 
    end process;
    type_cast_3146_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3146_inst_req_0;
      type_cast_3146_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3146_inst_req_1;
      type_cast_3146_inst_ack_1<= rack(0);
      type_cast_3146_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3146_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k840x_x0x_xph_3558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3146_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3150_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3150_inst_req_0;
      type_cast_3150_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3150_inst_req_1;
      type_cast_3150_inst_ack_1<= rack(0);
      type_cast_3150_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3150_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i844x_x1x_xph_3565,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3150_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3152_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3152_inst_req_0;
      type_cast_3152_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3152_inst_req_1;
      type_cast_3152_inst_ack_1<= rack(0);
      type_cast_3152_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3152_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div847_3023,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3152_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3156_inst_req_0;
      type_cast_3156_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3156_inst_req_1;
      type_cast_3156_inst_ack_1<= rack(0);
      type_cast_3156_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3156_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j894x_x0x_xph_3571,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3156_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3164_inst_req_0;
      type_cast_3164_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3164_inst_req_1;
      type_cast_3164_inst_ack_1<= rack(0);
      type_cast_3164_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3164_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3163_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv900_3165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3168_inst
    process(conv900_3165) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv900_3165(31 downto 0);
      type_cast_3168_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3170_inst
    process(conv902_3096) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv902_3096(31 downto 0);
      type_cast_3170_wire <= tmp_var; -- 
    end process;
    type_cast_3185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3185_inst_req_0;
      type_cast_3185_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3185_inst_req_1;
      type_cast_3185_inst_ack_1<= rack(0);
      type_cast_3185_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3185_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp908_3182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv909_3186,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3206_inst
    process(conv900_3165) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv900_3165(31 downto 0);
      type_cast_3206_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3208_inst
    process(add914_3203) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add914_3203(31 downto 0);
      type_cast_3208_wire <= tmp_var; -- 
    end process;
    type_cast_3221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3221_inst_req_0;
      type_cast_3221_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3221_inst_req_1;
      type_cast_3221_inst_ack_1<= rack(0);
      type_cast_3221_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3221_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3220_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv919_3222,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3225_inst
    process(conv919_3222) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv919_3222(31 downto 0);
      type_cast_3225_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3227_inst
    process(conv902_3096) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv902_3096(31 downto 0);
      type_cast_3227_wire <= tmp_var; -- 
    end process;
    type_cast_3242_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3242_inst_req_0;
      type_cast_3242_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3242_inst_req_1;
      type_cast_3242_inst_ack_1<= rack(0);
      type_cast_3242_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3242_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp927_3239,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv928_3243,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3257_inst
    process(conv919_3222) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv919_3222(31 downto 0);
      type_cast_3257_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3259_inst
    process(add932_3254) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add932_3254(31 downto 0);
      type_cast_3259_wire <= tmp_var; -- 
    end process;
    type_cast_3272_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3272_inst_req_0;
      type_cast_3272_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3272_inst_req_1;
      type_cast_3272_inst_ack_1<= rack(0);
      type_cast_3272_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3272_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3271_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv939_3273,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3277_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3277_inst_req_0;
      type_cast_3277_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3277_inst_req_1;
      type_cast_3277_inst_ack_1<= rack(0);
      type_cast_3277_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3277_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3276_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv943_3278,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3301_inst
    process(add951_3298) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add951_3298(31 downto 0);
      type_cast_3301_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3306_inst
    process(ASHR_i32_i32_3305_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3305_wire(31 downto 0);
      shr953_3307 <= tmp_var; -- 
    end process;
    type_cast_3311_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3311_inst_req_0;
      type_cast_3311_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3311_inst_req_1;
      type_cast_3311_inst_ack_1<= rack(0);
      type_cast_3311_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3311_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3310_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom954_3312,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3330_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3330_inst_req_0;
      type_cast_3330_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3330_inst_req_1;
      type_cast_3330_inst_ack_1<= rack(0);
      type_cast_3330_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3330_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3329_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv960_3331,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3384_inst
    process(add978_3361) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add978_3361(31 downto 0);
      type_cast_3384_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3389_inst
    process(ASHR_i32_i32_3388_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3388_wire(31 downto 0);
      shr996_3390 <= tmp_var; -- 
    end process;
    type_cast_3394_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3394_inst_req_0;
      type_cast_3394_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3394_inst_req_1;
      type_cast_3394_inst_ack_1<= rack(0);
      type_cast_3394_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3394_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3393_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom997_3395,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3409_inst
    process(add994_3381) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add994_3381(31 downto 0);
      type_cast_3409_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3414_inst
    process(ASHR_i32_i32_3413_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3413_wire(31 downto 0);
      shr1001_3415 <= tmp_var; -- 
    end process;
    type_cast_3419_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3419_inst_req_0;
      type_cast_3419_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3419_inst_req_1;
      type_cast_3419_inst_ack_1<= rack(0);
      type_cast_3419_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3419_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3418_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1002_3420,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3437_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3437_inst_req_0;
      type_cast_3437_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3437_inst_req_1;
      type_cast_3437_inst_ack_1<= rack(0);
      type_cast_3437_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3437_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3436_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1008_3438,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3447_inst
    process(add1009_3444) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1009_3444(31 downto 0);
      type_cast_3447_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3449_inst
    process(conv880_3057) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv880_3057(31 downto 0);
      type_cast_3449_wire <= tmp_var; -- 
    end process;
    type_cast_3476_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3476_inst_req_0;
      type_cast_3476_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3476_inst_req_1;
      type_cast_3476_inst_ack_1<= rack(0);
      type_cast_3476_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3476_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3475_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1023_3477,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3483_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3483_inst_req_0;
      type_cast_3483_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3483_inst_req_1;
      type_cast_3483_inst_ack_1<= rack(0);
      type_cast_3483_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3483_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1024_3480,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1025_3484,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3503_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3503_inst_req_0;
      type_cast_3503_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3503_inst_req_1;
      type_cast_3503_inst_ack_1<= rack(0);
      type_cast_3503_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3503_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1031_3500,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1036_3504,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3520_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3520_inst_req_0;
      type_cast_3520_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3520_inst_req_1;
      type_cast_3520_inst_ack_1<= rack(0);
      type_cast_3520_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3520_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3519_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1039_3521,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3527_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3527_inst_req_0;
      type_cast_3527_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3527_inst_req_1;
      type_cast_3527_inst_ack_1<= rack(0);
      type_cast_3527_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3527_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1040_3524,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1041_3528,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3561_inst_req_0;
      type_cast_3561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3561_inst_req_1;
      type_cast_3561_inst_ack_1<= rack(0);
      type_cast_3561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1017_3464,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3561_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3568_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3568_inst_req_0;
      type_cast_3568_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3568_inst_req_1;
      type_cast_3568_inst_ack_1<= rack(0);
      type_cast_3568_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3568_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i844x_x2_3147,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3568_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3570_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3570_inst_req_0;
      type_cast_3570_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3570_inst_req_1;
      type_cast_3570_inst_ack_1<= rack(0);
      type_cast_3570_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3570_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1036x_xi844x_x2_3509,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3570_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3574_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3574_inst_req_0;
      type_cast_3574_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3574_inst_req_1;
      type_cast_3574_inst_ack_1<= rack(0);
      type_cast_3574_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3574_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j894x_x2_3516,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3574_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3576_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3576_inst_req_0;
      type_cast_3576_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3576_inst_req_1;
      type_cast_3576_inst_ack_1<= rack(0);
      type_cast_3576_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3576_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j894x_x1_3153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3576_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3583_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3583_inst_req_0;
      type_cast_3583_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3583_inst_req_1;
      type_cast_3583_inst_ack_1<= rack(0);
      type_cast_3583_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3583_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1040_3524,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3583_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3587_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3587_inst_req_0;
      type_cast_3587_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3587_inst_req_1;
      type_cast_3587_inst_ack_1<= rack(0);
      type_cast_3587_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3587_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv1025_3484,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3587_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3591_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3591_inst_req_0;
      type_cast_3591_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3591_inst_req_1;
      type_cast_3591_inst_ack_1<= rack(0);
      type_cast_3591_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3591_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1024_3480,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3591_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3595_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3595_inst_req_0;
      type_cast_3595_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3595_inst_req_1;
      type_cast_3595_inst_ack_1<= rack(0);
      type_cast_3595_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3595_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1024x_xlcssa_3588,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1064_3596,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3605_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3605_inst_req_0;
      type_cast_3605_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3605_inst_req_1;
      type_cast_3605_inst_ack_1<= rack(0);
      type_cast_3605_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3605_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1040x_xlcssa_3580,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1070_3606,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3645_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3645_inst_req_0;
      type_cast_3645_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3645_inst_req_1;
      type_cast_3645_inst_ack_1<= rack(0);
      type_cast_3645_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3645_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1079_3618,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1104_3646,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3655_inst
    process(sext1774_3652) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1774_3652(31 downto 0);
      type_cast_3655_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3660_inst
    process(ASHR_i32_i32_3659_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3659_wire(31 downto 0);
      conv1112_3661 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3670_inst
    process(sext1726_3667) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1726_3667(31 downto 0);
      type_cast_3670_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3675_inst
    process(ASHR_i32_i32_3674_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3674_wire(31 downto 0);
      conv1114_3676 <= tmp_var; -- 
    end process;
    type_cast_3684_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3684_inst_req_0;
      type_cast_3684_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3684_inst_req_1;
      type_cast_3684_inst_ack_1<= rack(0);
      type_cast_3684_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3684_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1075_3615,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1126_3685,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3694_inst
    process(sext1775_3691) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1775_3691(31 downto 0);
      type_cast_3694_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3699_inst
    process(ASHR_i32_i32_3698_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3698_wire(31 downto 0);
      conv1170_3700 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3720_inst
    process(sext1727_3717) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1727_3717(31 downto 0);
      type_cast_3720_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3725_inst
    process(ASHR_i32_i32_3724_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3724_wire(31 downto 0);
      conv1194_3726 <= tmp_var; -- 
    end process;
    type_cast_3732_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3732_inst_req_0;
      type_cast_3732_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3732_inst_req_1;
      type_cast_3732_inst_ack_1<= rack(0);
      type_cast_3732_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3732_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k1060x_x0x_xph_4133,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3732_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3739_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3739_inst_req_0;
      type_cast_3739_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3739_inst_req_1;
      type_cast_3739_inst_ack_1<= rack(0);
      type_cast_3739_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3739_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1068x_x1x_xph_4140,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3739_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3741_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3741_inst_req_0;
      type_cast_3741_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3741_inst_req_1;
      type_cast_3741_inst_ack_1<= rack(0);
      type_cast_3741_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3741_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div1071_3612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3741_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3745_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3745_inst_req_0;
      type_cast_3745_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3745_inst_req_1;
      type_cast_3745_inst_ack_1<= rack(0);
      type_cast_3745_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3745_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div1065_3602,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3745_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3747_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3747_inst_req_0;
      type_cast_3747_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3747_inst_req_1;
      type_cast_3747_inst_ack_1<= rack(0);
      type_cast_3747_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3747_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1118x_x0x_xph_4146,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3747_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3752_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3752_inst_req_0;
      type_cast_3752_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3752_inst_req_1;
      type_cast_3752_inst_ack_1<= rack(0);
      type_cast_3752_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3752_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3751_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1124_3753,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3756_inst
    process(conv1124_3753) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1124_3753(31 downto 0);
      type_cast_3756_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3758_inst
    process(conv1126_3685) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1126_3685(31 downto 0);
      type_cast_3758_wire <= tmp_var; -- 
    end process;
    type_cast_3773_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3773_inst_req_0;
      type_cast_3773_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3773_inst_req_1;
      type_cast_3773_inst_ack_1<= rack(0);
      type_cast_3773_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3773_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1132_3770,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1133_3774,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3794_inst
    process(conv1124_3753) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1124_3753(31 downto 0);
      type_cast_3794_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3796_inst
    process(add1138_3791) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1138_3791(31 downto 0);
      type_cast_3796_wire <= tmp_var; -- 
    end process;
    type_cast_3809_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3809_inst_req_0;
      type_cast_3809_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3809_inst_req_1;
      type_cast_3809_inst_ack_1<= rack(0);
      type_cast_3809_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3809_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3808_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1143_3810,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3813_inst
    process(conv1143_3810) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1143_3810(31 downto 0);
      type_cast_3813_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3815_inst
    process(conv1126_3685) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1126_3685(31 downto 0);
      type_cast_3815_wire <= tmp_var; -- 
    end process;
    type_cast_3830_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3830_inst_req_0;
      type_cast_3830_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3830_inst_req_1;
      type_cast_3830_inst_ack_1<= rack(0);
      type_cast_3830_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3830_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1151_3827,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1152_3831,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3839_inst
    process(conv1143_3810) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1143_3810(31 downto 0);
      type_cast_3839_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3841_inst
    process(add1155_3836) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1155_3836(31 downto 0);
      type_cast_3841_wire <= tmp_var; -- 
    end process;
    type_cast_3854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3854_inst_req_0;
      type_cast_3854_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3854_inst_req_1;
      type_cast_3854_inst_ack_1<= rack(0);
      type_cast_3854_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3854_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3853_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1162_3855,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3859_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3859_inst_req_0;
      type_cast_3859_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3859_inst_req_1;
      type_cast_3859_inst_ack_1<= rack(0);
      type_cast_3859_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3859_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3858_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1166_3860,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3883_inst
    process(add1174_3880) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1174_3880(31 downto 0);
      type_cast_3883_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3888_inst
    process(ASHR_i32_i32_3887_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3887_wire(31 downto 0);
      shr1176_3889 <= tmp_var; -- 
    end process;
    type_cast_3893_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3893_inst_req_0;
      type_cast_3893_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3893_inst_req_1;
      type_cast_3893_inst_ack_1<= rack(0);
      type_cast_3893_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3893_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3892_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1177_3894,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3912_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3912_inst_req_0;
      type_cast_3912_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3912_inst_req_1;
      type_cast_3912_inst_ack_1<= rack(0);
      type_cast_3912_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3912_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3911_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1183_3913,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3966_inst
    process(add1201_3943) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1201_3943(31 downto 0);
      type_cast_3966_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3971_inst
    process(ASHR_i32_i32_3970_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3970_wire(31 downto 0);
      shr1219_3972 <= tmp_var; -- 
    end process;
    type_cast_3976_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3976_inst_req_0;
      type_cast_3976_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3976_inst_req_1;
      type_cast_3976_inst_ack_1<= rack(0);
      type_cast_3976_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3976_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3975_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1220_3977,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3991_inst
    process(add1217_3963) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1217_3963(31 downto 0);
      type_cast_3991_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3996_inst
    process(ASHR_i32_i32_3995_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3995_wire(31 downto 0);
      shr1224_3997 <= tmp_var; -- 
    end process;
    type_cast_4001_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4001_inst_req_0;
      type_cast_4001_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4001_inst_req_1;
      type_cast_4001_inst_ack_1<= rack(0);
      type_cast_4001_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4001_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4000_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1225_4002,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4019_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4019_inst_req_0;
      type_cast_4019_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4019_inst_req_1;
      type_cast_4019_inst_ack_1<= rack(0);
      type_cast_4019_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4019_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4018_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1231_4020,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4029_inst
    process(add1232_4026) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1232_4026(31 downto 0);
      type_cast_4029_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4031_inst
    process(conv1104_3646) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1104_3646(31 downto 0);
      type_cast_4031_wire <= tmp_var; -- 
    end process;
    type_cast_4058_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4058_inst_req_0;
      type_cast_4058_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4058_inst_req_1;
      type_cast_4058_inst_ack_1<= rack(0);
      type_cast_4058_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4058_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4057_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1246_4059,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4065_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4065_inst_req_0;
      type_cast_4065_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4065_inst_req_1;
      type_cast_4065_inst_ack_1<= rack(0);
      type_cast_4065_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4065_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1247_4062,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1248_4066,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4079_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4079_inst_req_0;
      type_cast_4079_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4079_inst_req_1;
      type_cast_4079_inst_ack_1<= rack(0);
      type_cast_4079_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4079_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1253_4076,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1258_4080,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4095_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4095_inst_req_0;
      type_cast_4095_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4095_inst_req_1;
      type_cast_4095_inst_ack_1<= rack(0);
      type_cast_4095_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4095_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4094_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1261_4096,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4102_inst_req_0;
      type_cast_4102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4102_inst_req_1;
      type_cast_4102_inst_ack_1<= rack(0);
      type_cast_4102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1262_4099,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1263_4103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4136_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4136_inst_req_0;
      type_cast_4136_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4136_inst_req_1;
      type_cast_4136_inst_ack_1<= rack(0);
      type_cast_4136_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4136_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1240_4046,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4136_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4143_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4143_inst_req_0;
      type_cast_4143_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4143_inst_req_1;
      type_cast_4143_inst_ack_1<= rack(0);
      type_cast_4143_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4143_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1068x_x2_3736,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4143_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4145_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4145_inst_req_0;
      type_cast_4145_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4145_inst_req_1;
      type_cast_4145_inst_ack_1<= rack(0);
      type_cast_4145_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4145_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1258x_xi1068x_x2_4085,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4145_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4149_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4149_inst_req_0;
      type_cast_4149_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4149_inst_req_1;
      type_cast_4149_inst_ack_1<= rack(0);
      type_cast_4149_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4149_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1118x_x1_3742,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4149_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4151_inst_req_0;
      type_cast_4151_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4151_inst_req_1;
      type_cast_4151_inst_ack_1<= rack(0);
      type_cast_4151_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4151_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1118x_x2_4091,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4151_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4158_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4158_inst_req_0;
      type_cast_4158_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4158_inst_req_1;
      type_cast_4158_inst_ack_1<= rack(0);
      type_cast_4158_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4158_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1262_4099,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4158_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4162_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4162_inst_req_0;
      type_cast_4162_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4162_inst_req_1;
      type_cast_4162_inst_ack_1<= rack(0);
      type_cast_4162_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4162_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv1248_4066,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4162_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4166_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4166_inst_req_0;
      type_cast_4166_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4166_inst_req_1;
      type_cast_4166_inst_ack_1<= rack(0);
      type_cast_4166_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4166_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1262x_xlcssa_4155,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1288_4167,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4212_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4212_inst_req_0;
      type_cast_4212_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4212_inst_req_1;
      type_cast_4212_inst_ack_1<= rack(0);
      type_cast_4212_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4212_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1298_4185,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1323_4213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4222_inst
    process(sext1776_4219) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1776_4219(31 downto 0);
      type_cast_4222_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4227_inst
    process(ASHR_i32_i32_4226_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4226_wire(31 downto 0);
      conv1331_4228 <= tmp_var; -- 
    end process;
    -- interlock type_cast_4237_inst
    process(sext1728_4234) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1728_4234(31 downto 0);
      type_cast_4237_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4242_inst
    process(ASHR_i32_i32_4241_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4241_wire(31 downto 0);
      conv1333_4243 <= tmp_var; -- 
    end process;
    type_cast_4251_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4251_inst_req_0;
      type_cast_4251_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4251_inst_req_1;
      type_cast_4251_inst_ack_1<= rack(0);
      type_cast_4251_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4251_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1294_4182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1345_4252,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4261_inst
    process(sext1777_4258) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1777_4258(31 downto 0);
      type_cast_4261_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4266_inst
    process(ASHR_i32_i32_4265_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4265_wire(31 downto 0);
      conv1388_4267 <= tmp_var; -- 
    end process;
    -- interlock type_cast_4287_inst
    process(sext1729_4284) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1729_4284(31 downto 0);
      type_cast_4287_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4292_inst
    process(ASHR_i32_i32_4291_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4291_wire(31 downto 0);
      conv1412_4293 <= tmp_var; -- 
    end process;
    type_cast_4302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4302_inst_req_0;
      type_cast_4302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4302_inst_req_1;
      type_cast_4302_inst_ack_1<= rack(0);
      type_cast_4302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k1282x_x0x_xph_4690,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4302_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4306_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4306_inst_req_0;
      type_cast_4306_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4306_inst_req_1;
      type_cast_4306_inst_ack_1<= rack(0);
      type_cast_4306_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4306_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul1290_4179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4306_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4308_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4308_inst_req_0;
      type_cast_4308_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4308_inst_req_1;
      type_cast_4308_inst_ack_1<= rack(0);
      type_cast_4308_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4308_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1286x_x1x_xph_4697,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4308_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4315_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4315_inst_req_0;
      type_cast_4315_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4315_inst_req_1;
      type_cast_4315_inst_ack_1<= rack(0);
      type_cast_4315_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4315_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1337x_x0x_xph_4703,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4315_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4320_inst_req_0;
      type_cast_4320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4320_inst_req_1;
      type_cast_4320_inst_ack_1<= rack(0);
      type_cast_4320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4319_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1343_4321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4324_inst
    process(conv1343_4321) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1343_4321(31 downto 0);
      type_cast_4324_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4326_inst
    process(conv1345_4252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1345_4252(31 downto 0);
      type_cast_4326_wire <= tmp_var; -- 
    end process;
    type_cast_4341_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4341_inst_req_0;
      type_cast_4341_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4341_inst_req_1;
      type_cast_4341_inst_ack_1<= rack(0);
      type_cast_4341_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4341_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1351_4338,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1352_4342,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4350_inst
    process(conv1343_4321) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1343_4321(31 downto 0);
      type_cast_4350_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4352_inst
    process(add1355_4347) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1355_4347(31 downto 0);
      type_cast_4352_wire <= tmp_var; -- 
    end process;
    type_cast_4365_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4365_inst_req_0;
      type_cast_4365_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4365_inst_req_1;
      type_cast_4365_inst_ack_1<= rack(0);
      type_cast_4365_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4365_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4364_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1360_4366,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4369_inst
    process(conv1360_4366) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1360_4366(31 downto 0);
      type_cast_4369_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4371_inst
    process(conv1345_4252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1345_4252(31 downto 0);
      type_cast_4371_wire <= tmp_var; -- 
    end process;
    type_cast_4386_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4386_inst_req_0;
      type_cast_4386_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4386_inst_req_1;
      type_cast_4386_inst_ack_1<= rack(0);
      type_cast_4386_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4386_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1368_4383,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1369_4387,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4401_inst
    process(conv1360_4366) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1360_4366(31 downto 0);
      type_cast_4401_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4403_inst
    process(add1373_4398) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1373_4398(31 downto 0);
      type_cast_4403_wire <= tmp_var; -- 
    end process;
    type_cast_4416_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4416_inst_req_0;
      type_cast_4416_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4416_inst_req_1;
      type_cast_4416_inst_ack_1<= rack(0);
      type_cast_4416_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4416_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4415_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1380_4417,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4421_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4421_inst_req_0;
      type_cast_4421_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4421_inst_req_1;
      type_cast_4421_inst_ack_1<= rack(0);
      type_cast_4421_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4421_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4420_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1384_4422,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4445_inst
    process(add1392_4442) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1392_4442(31 downto 0);
      type_cast_4445_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4450_inst
    process(ASHR_i32_i32_4449_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4449_wire(31 downto 0);
      shr1394_4451 <= tmp_var; -- 
    end process;
    type_cast_4455_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4455_inst_req_0;
      type_cast_4455_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4455_inst_req_1;
      type_cast_4455_inst_ack_1<= rack(0);
      type_cast_4455_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4455_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4454_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1395_4456,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4474_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4474_inst_req_0;
      type_cast_4474_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4474_inst_req_1;
      type_cast_4474_inst_ack_1<= rack(0);
      type_cast_4474_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4474_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4473_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1401_4475,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4528_inst
    process(add1419_4505) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1419_4505(31 downto 0);
      type_cast_4528_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4533_inst
    process(ASHR_i32_i32_4532_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4532_wire(31 downto 0);
      shr1437_4534 <= tmp_var; -- 
    end process;
    type_cast_4538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4538_inst_req_0;
      type_cast_4538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4538_inst_req_1;
      type_cast_4538_inst_ack_1<= rack(0);
      type_cast_4538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4537_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1438_4539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4553_inst
    process(add1435_4525) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1435_4525(31 downto 0);
      type_cast_4553_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4558_inst
    process(ASHR_i32_i32_4557_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4557_wire(31 downto 0);
      shr1442_4559 <= tmp_var; -- 
    end process;
    type_cast_4563_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4563_inst_req_0;
      type_cast_4563_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4563_inst_req_1;
      type_cast_4563_inst_ack_1<= rack(0);
      type_cast_4563_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4563_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4562_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1443_4564,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4581_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4581_inst_req_0;
      type_cast_4581_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4581_inst_req_1;
      type_cast_4581_inst_ack_1<= rack(0);
      type_cast_4581_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4581_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4580_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1449_4582,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4591_inst
    process(add1450_4588) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1450_4588(31 downto 0);
      type_cast_4591_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4593_inst
    process(conv1323_4213) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1323_4213(31 downto 0);
      type_cast_4593_wire <= tmp_var; -- 
    end process;
    type_cast_4620_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4620_inst_req_0;
      type_cast_4620_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4620_inst_req_1;
      type_cast_4620_inst_ack_1<= rack(0);
      type_cast_4620_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4620_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4619_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1464_4621,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4627_inst_req_0;
      type_cast_4627_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4627_inst_req_1;
      type_cast_4627_inst_ack_1<= rack(0);
      type_cast_4627_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4627_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1465_4624,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1466_4628,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4647_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4647_inst_req_0;
      type_cast_4647_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4647_inst_req_1;
      type_cast_4647_inst_ack_1<= rack(0);
      type_cast_4647_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4647_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1472_4644,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1477_4648,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4664_inst_req_0;
      type_cast_4664_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4664_inst_req_1;
      type_cast_4664_inst_ack_1<= rack(0);
      type_cast_4664_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4664_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4663_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1480_4665,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4671_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4671_inst_req_0;
      type_cast_4671_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4671_inst_req_1;
      type_cast_4671_inst_ack_1<= rack(0);
      type_cast_4671_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4671_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1481_4668,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1482_4672,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4696_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4696_inst_req_0;
      type_cast_4696_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4696_inst_req_1;
      type_cast_4696_inst_ack_1<= rack(0);
      type_cast_4696_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4696_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1458_4608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4696_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4700_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4700_inst_req_0;
      type_cast_4700_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4700_inst_req_1;
      type_cast_4700_inst_ack_1<= rack(0);
      type_cast_4700_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4700_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1286x_x2_4303,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4700_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4702_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4702_inst_req_0;
      type_cast_4702_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4702_inst_req_1;
      type_cast_4702_inst_ack_1<= rack(0);
      type_cast_4702_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4702_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1477x_xi1286x_x2_4653,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4702_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4706_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4706_inst_req_0;
      type_cast_4706_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4706_inst_req_1;
      type_cast_4706_inst_ack_1<= rack(0);
      type_cast_4706_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4706_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1337x_x2_4660,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4706_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4708_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4708_inst_req_0;
      type_cast_4708_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4708_inst_req_1;
      type_cast_4708_inst_ack_1<= rack(0);
      type_cast_4708_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4708_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1337x_x1_4309,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4708_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4715_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4715_inst_req_0;
      type_cast_4715_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4715_inst_req_1;
      type_cast_4715_inst_ack_1<= rack(0);
      type_cast_4715_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4715_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1481_4668,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4715_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4719_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4719_inst_req_0;
      type_cast_4719_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4719_inst_req_1;
      type_cast_4719_inst_ack_1<= rack(0);
      type_cast_4719_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4719_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv1466_4628,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4719_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4723_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4723_inst_req_0;
      type_cast_4723_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4723_inst_req_1;
      type_cast_4723_inst_ack_1<= rack(0);
      type_cast_4723_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4723_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1465_4624,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4723_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4727_inst_req_0;
      type_cast_4727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4727_inst_req_1;
      type_cast_4727_inst_ack_1<= rack(0);
      type_cast_4727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1465x_xlcssa_4720,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1503_4728,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4737_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4737_inst_req_0;
      type_cast_4737_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4737_inst_req_1;
      type_cast_4737_inst_ack_1<= rack(0);
      type_cast_4737_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4737_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1481x_xlcssa_4712,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1509_4738,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4783_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4783_inst_req_0;
      type_cast_4783_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4783_inst_req_1;
      type_cast_4783_inst_ack_1<= rack(0);
      type_cast_4783_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4783_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1519_4756,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1544_4784,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4793_inst
    process(sext1778_4790) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1778_4790(31 downto 0);
      type_cast_4793_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4798_inst
    process(ASHR_i32_i32_4797_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4797_wire(31 downto 0);
      conv1552_4799 <= tmp_var; -- 
    end process;
    -- interlock type_cast_4808_inst
    process(sext1730_4805) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1730_4805(31 downto 0);
      type_cast_4808_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4813_inst
    process(ASHR_i32_i32_4812_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4812_wire(31 downto 0);
      conv1554_4814 <= tmp_var; -- 
    end process;
    type_cast_4822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4822_inst_req_0;
      type_cast_4822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4822_inst_req_1;
      type_cast_4822_inst_ack_1<= rack(0);
      type_cast_4822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4822_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1515_4753,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1566_4823,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4832_inst
    process(sext1779_4829) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1779_4829(31 downto 0);
      type_cast_4832_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4837_inst
    process(ASHR_i32_i32_4836_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4836_wire(31 downto 0);
      conv1608_4838 <= tmp_var; -- 
    end process;
    -- interlock type_cast_4858_inst
    process(sext1731_4855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1731_4855(31 downto 0);
      type_cast_4858_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4863_inst
    process(ASHR_i32_i32_4862_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4862_wire(31 downto 0);
      conv1632_4864 <= tmp_var; -- 
    end process;
    type_cast_4873_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4873_inst_req_0;
      type_cast_4873_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4873_inst_req_1;
      type_cast_4873_inst_ack_1<= rack(0);
      type_cast_4873_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4873_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k1499x_x0x_xph_5247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4873_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4877_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4877_inst_req_0;
      type_cast_4877_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4877_inst_req_1;
      type_cast_4877_inst_ack_1<= rack(0);
      type_cast_4877_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4877_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div1511_4750,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4877_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4879_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4879_inst_req_0;
      type_cast_4879_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4879_inst_req_1;
      type_cast_4879_inst_ack_1<= rack(0);
      type_cast_4879_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4879_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1507x_x1x_xph_5254,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4879_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4883_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4883_inst_req_0;
      type_cast_4883_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4883_inst_req_1;
      type_cast_4883_inst_ack_1<= rack(0);
      type_cast_4883_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4883_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1558x_x0x_xph_5260,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4883_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4885_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4885_inst_req_0;
      type_cast_4885_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4885_inst_req_1;
      type_cast_4885_inst_ack_1<= rack(0);
      type_cast_4885_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4885_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div1504_4734,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4885_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4890_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4890_inst_req_0;
      type_cast_4890_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4890_inst_req_1;
      type_cast_4890_inst_ack_1<= rack(0);
      type_cast_4890_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4890_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4889_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1564_4891,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4894_inst
    process(conv1564_4891) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1564_4891(31 downto 0);
      type_cast_4894_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4896_inst
    process(conv1566_4823) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1566_4823(31 downto 0);
      type_cast_4896_wire <= tmp_var; -- 
    end process;
    type_cast_4911_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4911_inst_req_0;
      type_cast_4911_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4911_inst_req_1;
      type_cast_4911_inst_ack_1<= rack(0);
      type_cast_4911_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4911_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1572_4908,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1573_4912,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4920_inst
    process(conv1564_4891) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1564_4891(31 downto 0);
      type_cast_4920_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4922_inst
    process(add1576_4917) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1576_4917(31 downto 0);
      type_cast_4922_wire <= tmp_var; -- 
    end process;
    type_cast_4935_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4935_inst_req_0;
      type_cast_4935_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4935_inst_req_1;
      type_cast_4935_inst_ack_1<= rack(0);
      type_cast_4935_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4935_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4934_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1581_4936,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4939_inst
    process(conv1581_4936) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1581_4936(31 downto 0);
      type_cast_4939_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4941_inst
    process(conv1566_4823) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1566_4823(31 downto 0);
      type_cast_4941_wire <= tmp_var; -- 
    end process;
    type_cast_4956_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4956_inst_req_0;
      type_cast_4956_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4956_inst_req_1;
      type_cast_4956_inst_ack_1<= rack(0);
      type_cast_4956_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4956_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1589_4953,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1590_4957,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4965_inst
    process(conv1581_4936) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1581_4936(31 downto 0);
      type_cast_4965_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4967_inst
    process(add1593_4962) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1593_4962(31 downto 0);
      type_cast_4967_wire <= tmp_var; -- 
    end process;
    type_cast_4980_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4980_inst_req_0;
      type_cast_4980_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4980_inst_req_1;
      type_cast_4980_inst_ack_1<= rack(0);
      type_cast_4980_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4980_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4979_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1600_4981,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4985_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4985_inst_req_0;
      type_cast_4985_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4985_inst_req_1;
      type_cast_4985_inst_ack_1<= rack(0);
      type_cast_4985_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4985_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4984_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1604_4986,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_5009_inst
    process(add1612_5006) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1612_5006(31 downto 0);
      type_cast_5009_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_5014_inst
    process(ASHR_i32_i32_5013_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_5013_wire(31 downto 0);
      shr1614_5015 <= tmp_var; -- 
    end process;
    type_cast_5019_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5019_inst_req_0;
      type_cast_5019_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5019_inst_req_1;
      type_cast_5019_inst_ack_1<= rack(0);
      type_cast_5019_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5019_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5018_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1615_5020,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5038_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5038_inst_req_0;
      type_cast_5038_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5038_inst_req_1;
      type_cast_5038_inst_ack_1<= rack(0);
      type_cast_5038_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5038_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5037_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1621_5039,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_5092_inst
    process(add1639_5069) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1639_5069(31 downto 0);
      type_cast_5092_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_5097_inst
    process(ASHR_i32_i32_5096_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_5096_wire(31 downto 0);
      shr1657_5098 <= tmp_var; -- 
    end process;
    type_cast_5102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5102_inst_req_0;
      type_cast_5102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5102_inst_req_1;
      type_cast_5102_inst_ack_1<= rack(0);
      type_cast_5102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5101_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1658_5103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_5117_inst
    process(add1655_5089) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1655_5089(31 downto 0);
      type_cast_5117_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_5122_inst
    process(ASHR_i32_i32_5121_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_5121_wire(31 downto 0);
      shr1662_5123 <= tmp_var; -- 
    end process;
    type_cast_5127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5127_inst_req_0;
      type_cast_5127_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5127_inst_req_1;
      type_cast_5127_inst_ack_1<= rack(0);
      type_cast_5127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5126_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1663_5128,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5145_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5145_inst_req_0;
      type_cast_5145_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5145_inst_req_1;
      type_cast_5145_inst_ack_1<= rack(0);
      type_cast_5145_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5145_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5144_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1669_5146,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_5155_inst
    process(add1670_5152) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1670_5152(31 downto 0);
      type_cast_5155_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_5157_inst
    process(conv1544_4784) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1544_4784(31 downto 0);
      type_cast_5157_wire <= tmp_var; -- 
    end process;
    type_cast_5184_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5184_inst_req_0;
      type_cast_5184_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5184_inst_req_1;
      type_cast_5184_inst_ack_1<= rack(0);
      type_cast_5184_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5184_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5183_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1684_5185,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5191_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5191_inst_req_0;
      type_cast_5191_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5191_inst_req_1;
      type_cast_5191_inst_ack_1<= rack(0);
      type_cast_5191_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5191_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1685_5188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1686_5192,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5205_inst_req_0;
      type_cast_5205_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5205_inst_req_1;
      type_cast_5205_inst_ack_1<= rack(0);
      type_cast_5205_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5205_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1691_5202,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1696_5206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5221_inst_req_0;
      type_cast_5221_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5221_inst_req_1;
      type_cast_5221_inst_ack_1<= rack(0);
      type_cast_5221_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5221_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5220_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1699_5222,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5228_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5228_inst_req_0;
      type_cast_5228_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5228_inst_req_1;
      type_cast_5228_inst_ack_1<= rack(0);
      type_cast_5228_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5228_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1700_5225,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1701_5229,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5250_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5250_inst_req_0;
      type_cast_5250_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5250_inst_req_1;
      type_cast_5250_inst_ack_1<= rack(0);
      type_cast_5250_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5250_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1678_5172,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_5250_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5257_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5257_inst_req_0;
      type_cast_5257_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5257_inst_req_1;
      type_cast_5257_inst_ack_1<= rack(0);
      type_cast_5257_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5257_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1507x_x2_4874,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_5257_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5259_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5259_inst_req_0;
      type_cast_5259_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5259_inst_req_1;
      type_cast_5259_inst_ack_1<= rack(0);
      type_cast_5259_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5259_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1696x_xi1507x_x2_5211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_5259_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5263_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5263_inst_req_0;
      type_cast_5263_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5263_inst_req_1;
      type_cast_5263_inst_ack_1<= rack(0);
      type_cast_5263_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5263_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1558x_x2_5217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_5263_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5265_inst_req_0;
      type_cast_5265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5265_inst_req_1;
      type_cast_5265_inst_ack_1<= rack(0);
      type_cast_5265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1558x_x1_4880,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_5265_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_731_inst_req_0;
      type_cast_731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_731_inst_req_1;
      type_cast_731_inst_ack_1<= rack(0);
      type_cast_731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_731_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_728,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_732,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_750_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_750_inst_req_0;
      type_cast_750_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_750_inst_req_1;
      type_cast_750_inst_ack_1<= rack(0);
      type_cast_750_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_750_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_747,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_751,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_769_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_769_inst_req_0;
      type_cast_769_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_769_inst_req_1;
      type_cast_769_inst_ack_1<= rack(0);
      type_cast_769_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_769_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_766,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_770,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_810_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_810_inst_req_0;
      type_cast_810_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_810_inst_req_1;
      type_cast_810_inst_ack_1<= rack(0);
      type_cast_810_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_810_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_780,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_811,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_814_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_814_inst_req_0;
      type_cast_814_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_814_inst_req_1;
      type_cast_814_inst_ack_1<= rack(0);
      type_cast_814_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_814_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp15_783,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_815,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_825_inst
    process(sext1764_821) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1764_821(31 downto 0);
      type_cast_825_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_830_inst
    process(ASHR_i32_i32_829_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_829_wire(31 downto 0);
      conv37_831 <= tmp_var; -- 
    end process;
    -- interlock type_cast_840_inst
    process(sext_837) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_837(31 downto 0);
      type_cast_840_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_845_inst
    process(ASHR_i32_i32_844_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_844_wire(31 downto 0);
      conv39_846 <= tmp_var; -- 
    end process;
    type_cast_854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_854_inst_req_0;
      type_cast_854_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_854_inst_req_1;
      type_cast_854_inst_ack_1<= rack(0);
      type_cast_854_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_854_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp9_777,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_855,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_864_inst
    process(sext1765_861) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1765_861(31 downto 0);
      type_cast_864_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_869_inst
    process(ASHR_i32_i32_868_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_868_wire(31 downto 0);
      conv86_870 <= tmp_var; -- 
    end process;
    -- interlock type_cast_890_inst
    process(sext1717_887) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1717_887(31 downto 0);
      type_cast_890_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_895_inst
    process(ASHR_i32_i32_894_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_894_wire(31 downto 0);
      conv104_896 <= tmp_var; -- 
    end process;
    type_cast_905_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_905_inst_req_0;
      type_cast_905_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_905_inst_req_1;
      type_cast_905_inst_ack_1<= rack(0);
      type_cast_905_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_905_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_1307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_905_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_912_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_912_inst_req_0;
      type_cast_912_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_912_inst_req_1;
      type_cast_912_inst_ack_1<= rack(0);
      type_cast_912_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_912_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_1313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_912_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_919_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_919_inst_req_0;
      type_cast_919_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_919_inst_req_1;
      type_cast_919_inst_ack_1<= rack(0);
      type_cast_919_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_919_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_1319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_919_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_924_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_924_inst_req_0;
      type_cast_924_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_924_inst_req_1;
      type_cast_924_inst_ack_1<= rack(0);
      type_cast_924_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_924_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_923_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv46_925,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_928_inst
    process(conv46_925) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv46_925(31 downto 0);
      type_cast_928_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_930_inst
    process(conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv48_855(31 downto 0);
      type_cast_930_wire <= tmp_var; -- 
    end process;
    type_cast_945_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_945_inst_req_0;
      type_cast_945_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_945_inst_req_1;
      type_cast_945_inst_ack_1<= rack(0);
      type_cast_945_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_945_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp52_942,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_946,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_960_inst
    process(conv46_925) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv46_925(31 downto 0);
      type_cast_960_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_962_inst
    process(add_957) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_957(31 downto 0);
      type_cast_962_wire <= tmp_var; -- 
    end process;
    type_cast_975_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_975_inst_req_0;
      type_cast_975_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_975_inst_req_1;
      type_cast_975_inst_ack_1<= rack(0);
      type_cast_975_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_975_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_974_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_976,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_979_inst
    process(conv60_976) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv60_976(31 downto 0);
      type_cast_979_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_981_inst
    process(conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv48_855(31 downto 0);
      type_cast_981_wire <= tmp_var; -- 
    end process;
    type_cast_996_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_996_inst_req_0;
      type_cast_996_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_996_inst_req_1;
      type_cast_996_inst_ack_1<= rack(0);
      type_cast_996_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_996_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp68_993,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_997,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_col_high_1234_gather_scatter
    process(LOAD_col_high_1234_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_1234_data_0;
      ov(7 downto 0) := iv;
      tmp154_1235 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_1556_gather_scatter
    process(LOAD_col_high_1556_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_1556_data_0;
      ov(7 downto 0) := iv;
      tmp272_1557 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_1791_gather_scatter
    process(LOAD_col_high_1791_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_1791_data_0;
      ov(7 downto 0) := iv;
      tmp368_1792 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_2106_gather_scatter
    process(LOAD_col_high_2106_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_2106_data_0;
      ov(7 downto 0) := iv;
      tmp488_2107 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_2347_gather_scatter
    process(LOAD_col_high_2347_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_2347_data_0;
      ov(7 downto 0) := iv;
      tmp585_2348 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_2682_gather_scatter
    process(LOAD_col_high_2682_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_2682_data_0;
      ov(7 downto 0) := iv;
      tmp710_2683 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_2917_gather_scatter
    process(LOAD_col_high_2917_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_2917_data_0;
      ov(7 downto 0) := iv;
      tmp806_2918 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_3238_gather_scatter
    process(LOAD_col_high_3238_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_3238_data_0;
      ov(7 downto 0) := iv;
      tmp927_3239 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_3479_gather_scatter
    process(LOAD_col_high_3479_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_3479_data_0;
      ov(7 downto 0) := iv;
      tmp1024_3480 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_3826_gather_scatter
    process(LOAD_col_high_3826_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_3826_data_0;
      ov(7 downto 0) := iv;
      tmp1151_3827 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4061_gather_scatter
    process(LOAD_col_high_4061_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4061_data_0;
      ov(7 downto 0) := iv;
      tmp1247_4062 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4382_gather_scatter
    process(LOAD_col_high_4382_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4382_data_0;
      ov(7 downto 0) := iv;
      tmp1368_4383 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4623_gather_scatter
    process(LOAD_col_high_4623_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4623_data_0;
      ov(7 downto 0) := iv;
      tmp1465_4624 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4952_gather_scatter
    process(LOAD_col_high_4952_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4952_data_0;
      ov(7 downto 0) := iv;
      tmp1589_4953 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_5187_gather_scatter
    process(LOAD_col_high_5187_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_5187_data_0;
      ov(7 downto 0) := iv;
      tmp1685_5188 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_782_gather_scatter
    process(LOAD_col_high_782_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_782_data_0;
      ov(7 downto 0) := iv;
      tmp15_783 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_992_gather_scatter
    process(LOAD_col_high_992_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_992_data_0;
      ov(7 downto 0) := iv;
      tmp68_993 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_1352_gather_scatter
    process(LOAD_depth_high_1352_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_1352_data_0;
      ov(7 downto 0) := iv;
      tmp201_1353 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_1902_gather_scatter
    process(LOAD_depth_high_1902_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_1902_data_0;
      ov(7 downto 0) := iv;
      tmp417_1903 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_2479_gather_scatter
    process(LOAD_depth_high_2479_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_2479_data_0;
      ov(7 downto 0) := iv;
      tmp639_2480 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_3028_gather_scatter
    process(LOAD_depth_high_3028_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_3028_data_0;
      ov(7 downto 0) := iv;
      tmp855_3029 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_3617_gather_scatter
    process(LOAD_depth_high_3617_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_3617_data_0;
      ov(7 downto 0) := iv;
      tmp1079_3618 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_4184_gather_scatter
    process(LOAD_depth_high_4184_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_4184_data_0;
      ov(7 downto 0) := iv;
      tmp1298_4185 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_4755_gather_scatter
    process(LOAD_depth_high_4755_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_4755_data_0;
      ov(7 downto 0) := iv;
      tmp1519_4756 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_779_gather_scatter
    process(LOAD_depth_high_779_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_779_data_0;
      ov(7 downto 0) := iv;
      tmp12_780 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_1349_gather_scatter
    process(LOAD_pad_1349_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_1349_data_0;
      ov(7 downto 0) := iv;
      tmp197_1350 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_1899_gather_scatter
    process(LOAD_pad_1899_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_1899_data_0;
      ov(7 downto 0) := iv;
      tmp413_1900 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_2476_gather_scatter
    process(LOAD_pad_2476_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_2476_data_0;
      ov(7 downto 0) := iv;
      tmp635_2477 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_3025_gather_scatter
    process(LOAD_pad_3025_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_3025_data_0;
      ov(7 downto 0) := iv;
      tmp851_3026 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_3614_gather_scatter
    process(LOAD_pad_3614_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_3614_data_0;
      ov(7 downto 0) := iv;
      tmp1075_3615 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_4181_gather_scatter
    process(LOAD_pad_4181_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_4181_data_0;
      ov(7 downto 0) := iv;
      tmp1294_4182 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_4752_gather_scatter
    process(LOAD_pad_4752_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_4752_data_0;
      ov(7 downto 0) := iv;
      tmp1515_4753 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_776_gather_scatter
    process(LOAD_pad_776_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_776_data_0;
      ov(7 downto 0) := iv;
      tmp9_777 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_1278_gather_scatter
    process(LOAD_row_high_1278_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_1278_data_0;
      ov(7 downto 0) := iv;
      tmp169_1279 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_1505_gather_scatter
    process(LOAD_row_high_1505_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_1505_data_0;
      ov(7 downto 0) := iv;
      tmp254_1506 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_1828_gather_scatter
    process(LOAD_row_high_1828_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_1828_data_0;
      ov(7 downto 0) := iv;
      tmp383_1829 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_2055_gather_scatter
    process(LOAD_row_high_2055_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_2055_data_0;
      ov(7 downto 0) := iv;
      tmp470_2056 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_2391_gather_scatter
    process(LOAD_row_high_2391_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_2391_data_0;
      ov(7 downto 0) := iv;
      tmp601_2392 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_2631_gather_scatter
    process(LOAD_row_high_2631_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_2631_data_0;
      ov(7 downto 0) := iv;
      tmp692_2632 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_2954_gather_scatter
    process(LOAD_row_high_2954_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_2954_data_0;
      ov(7 downto 0) := iv;
      tmp821_2955 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_3181_gather_scatter
    process(LOAD_row_high_3181_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_3181_data_0;
      ov(7 downto 0) := iv;
      tmp908_3182 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_3523_gather_scatter
    process(LOAD_row_high_3523_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_3523_data_0;
      ov(7 downto 0) := iv;
      tmp1040_3524 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_3769_gather_scatter
    process(LOAD_row_high_3769_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_3769_data_0;
      ov(7 downto 0) := iv;
      tmp1132_3770 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_4098_gather_scatter
    process(LOAD_row_high_4098_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_4098_data_0;
      ov(7 downto 0) := iv;
      tmp1262_4099 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_4337_gather_scatter
    process(LOAD_row_high_4337_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_4337_data_0;
      ov(7 downto 0) := iv;
      tmp1351_4338 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_4667_gather_scatter
    process(LOAD_row_high_4667_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_4667_data_0;
      ov(7 downto 0) := iv;
      tmp1481_4668 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_4907_gather_scatter
    process(LOAD_row_high_4907_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_4907_data_0;
      ov(7 downto 0) := iv;
      tmp1572_4908 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_5224_gather_scatter
    process(LOAD_row_high_5224_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_5224_data_0;
      ov(7 downto 0) := iv;
      tmp1700_5225 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_941_gather_scatter
    process(LOAD_row_high_941_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_941_data_0;
      ov(7 downto 0) := iv;
      tmp52_942 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_col_high_752_gather_scatter
    process(conv2_751) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv2_751;
      ov(7 downto 0) := iv;
      STORE_col_high_752_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_depth_high_771_gather_scatter
    process(conv4_770) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv4_770;
      ov(7 downto 0) := iv;
      STORE_depth_high_771_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_row_high_733_gather_scatter
    process(conv_732) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_732;
      ov(7 downto 0) := iv;
      STORE_row_high_733_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1072_index_1_rename
    process(R_idxprom_1071_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1071_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1071_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1072_index_1_resize
    process(idxprom_1067) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1067;
      ov := iv(13 downto 0);
      R_idxprom_1071_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1072_root_address_inst
    process(array_obj_ref_1072_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1072_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1072_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1155_index_1_rename
    process(R_idxprom130_1154_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom130_1154_resized;
      ov(13 downto 0) := iv;
      R_idxprom130_1154_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1155_index_1_resize
    process(idxprom130_1150) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom130_1150;
      ov := iv(13 downto 0);
      R_idxprom130_1154_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1155_root_address_inst
    process(array_obj_ref_1155_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1155_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1155_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1180_index_1_rename
    process(R_idxprom135_1179_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom135_1179_resized;
      ov(13 downto 0) := iv;
      R_idxprom135_1179_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1180_index_1_resize
    process(idxprom135_1175) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom135_1175;
      ov := iv(13 downto 0);
      R_idxprom135_1179_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1180_root_address_inst
    process(array_obj_ref_1180_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1180_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1180_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1629_index_1_rename
    process(R_idxprom298_1628_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom298_1628_resized;
      ov(13 downto 0) := iv;
      R_idxprom298_1628_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1629_index_1_resize
    process(idxprom298_1624) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom298_1624;
      ov := iv(13 downto 0);
      R_idxprom298_1628_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1629_root_address_inst
    process(array_obj_ref_1629_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1629_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1629_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1712_index_1_rename
    process(R_idxprom341_1711_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom341_1711_resized;
      ov(13 downto 0) := iv;
      R_idxprom341_1711_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1712_index_1_resize
    process(idxprom341_1707) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom341_1707;
      ov := iv(13 downto 0);
      R_idxprom341_1711_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1712_root_address_inst
    process(array_obj_ref_1712_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1712_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1712_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1737_index_1_rename
    process(R_idxprom346_1736_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom346_1736_resized;
      ov(13 downto 0) := iv;
      R_idxprom346_1736_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1737_index_1_resize
    process(idxprom346_1732) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom346_1732;
      ov := iv(13 downto 0);
      R_idxprom346_1736_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1737_root_address_inst
    process(array_obj_ref_1737_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1737_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1737_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2185_index_1_rename
    process(R_idxprom515_2184_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom515_2184_resized;
      ov(13 downto 0) := iv;
      R_idxprom515_2184_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2185_index_1_resize
    process(idxprom515_2180) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom515_2180;
      ov := iv(13 downto 0);
      R_idxprom515_2184_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2185_root_address_inst
    process(array_obj_ref_2185_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2185_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2185_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2268_index_1_rename
    process(R_idxprom558_2267_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom558_2267_resized;
      ov(13 downto 0) := iv;
      R_idxprom558_2267_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2268_index_1_resize
    process(idxprom558_2263) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom558_2263;
      ov := iv(13 downto 0);
      R_idxprom558_2267_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2268_root_address_inst
    process(array_obj_ref_2268_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2268_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2268_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2293_index_1_rename
    process(R_idxprom563_2292_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom563_2292_resized;
      ov(13 downto 0) := iv;
      R_idxprom563_2292_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2293_index_1_resize
    process(idxprom563_2288) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom563_2288;
      ov := iv(13 downto 0);
      R_idxprom563_2292_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2293_root_address_inst
    process(array_obj_ref_2293_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2293_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2293_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2755_index_1_rename
    process(R_idxprom736_2754_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom736_2754_resized;
      ov(13 downto 0) := iv;
      R_idxprom736_2754_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2755_index_1_resize
    process(idxprom736_2750) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom736_2750;
      ov := iv(13 downto 0);
      R_idxprom736_2754_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2755_root_address_inst
    process(array_obj_ref_2755_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2755_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2755_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2838_index_1_rename
    process(R_idxprom779_2837_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom779_2837_resized;
      ov(13 downto 0) := iv;
      R_idxprom779_2837_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2838_index_1_resize
    process(idxprom779_2833) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom779_2833;
      ov := iv(13 downto 0);
      R_idxprom779_2837_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2838_root_address_inst
    process(array_obj_ref_2838_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2838_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2838_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2863_index_1_rename
    process(R_idxprom784_2862_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom784_2862_resized;
      ov(13 downto 0) := iv;
      R_idxprom784_2862_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2863_index_1_resize
    process(idxprom784_2858) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom784_2858;
      ov := iv(13 downto 0);
      R_idxprom784_2862_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2863_root_address_inst
    process(array_obj_ref_2863_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2863_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2863_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3317_index_1_rename
    process(R_idxprom954_3316_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom954_3316_resized;
      ov(13 downto 0) := iv;
      R_idxprom954_3316_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3317_index_1_resize
    process(idxprom954_3312) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom954_3312;
      ov := iv(13 downto 0);
      R_idxprom954_3316_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3317_root_address_inst
    process(array_obj_ref_3317_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3317_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3317_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3400_index_1_rename
    process(R_idxprom997_3399_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom997_3399_resized;
      ov(13 downto 0) := iv;
      R_idxprom997_3399_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3400_index_1_resize
    process(idxprom997_3395) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom997_3395;
      ov := iv(13 downto 0);
      R_idxprom997_3399_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3400_root_address_inst
    process(array_obj_ref_3400_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3400_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3400_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3425_index_1_rename
    process(R_idxprom1002_3424_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1002_3424_resized;
      ov(13 downto 0) := iv;
      R_idxprom1002_3424_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3425_index_1_resize
    process(idxprom1002_3420) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1002_3420;
      ov := iv(13 downto 0);
      R_idxprom1002_3424_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3425_root_address_inst
    process(array_obj_ref_3425_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3425_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3425_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3899_index_1_rename
    process(R_idxprom1177_3898_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1177_3898_resized;
      ov(13 downto 0) := iv;
      R_idxprom1177_3898_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3899_index_1_resize
    process(idxprom1177_3894) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1177_3894;
      ov := iv(13 downto 0);
      R_idxprom1177_3898_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3899_root_address_inst
    process(array_obj_ref_3899_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3899_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3899_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3982_index_1_rename
    process(R_idxprom1220_3981_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1220_3981_resized;
      ov(13 downto 0) := iv;
      R_idxprom1220_3981_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3982_index_1_resize
    process(idxprom1220_3977) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1220_3977;
      ov := iv(13 downto 0);
      R_idxprom1220_3981_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3982_root_address_inst
    process(array_obj_ref_3982_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3982_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3982_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4007_index_1_rename
    process(R_idxprom1225_4006_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1225_4006_resized;
      ov(13 downto 0) := iv;
      R_idxprom1225_4006_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4007_index_1_resize
    process(idxprom1225_4002) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1225_4002;
      ov := iv(13 downto 0);
      R_idxprom1225_4006_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4007_root_address_inst
    process(array_obj_ref_4007_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4007_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4007_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4461_index_1_rename
    process(R_idxprom1395_4460_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1395_4460_resized;
      ov(13 downto 0) := iv;
      R_idxprom1395_4460_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4461_index_1_resize
    process(idxprom1395_4456) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1395_4456;
      ov := iv(13 downto 0);
      R_idxprom1395_4460_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4461_root_address_inst
    process(array_obj_ref_4461_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4461_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4461_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4544_index_1_rename
    process(R_idxprom1438_4543_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1438_4543_resized;
      ov(13 downto 0) := iv;
      R_idxprom1438_4543_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4544_index_1_resize
    process(idxprom1438_4539) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1438_4539;
      ov := iv(13 downto 0);
      R_idxprom1438_4543_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4544_root_address_inst
    process(array_obj_ref_4544_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4544_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4544_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4569_index_1_rename
    process(R_idxprom1443_4568_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1443_4568_resized;
      ov(13 downto 0) := iv;
      R_idxprom1443_4568_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4569_index_1_resize
    process(idxprom1443_4564) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1443_4564;
      ov := iv(13 downto 0);
      R_idxprom1443_4568_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4569_root_address_inst
    process(array_obj_ref_4569_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4569_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4569_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5025_index_1_rename
    process(R_idxprom1615_5024_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1615_5024_resized;
      ov(13 downto 0) := iv;
      R_idxprom1615_5024_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5025_index_1_resize
    process(idxprom1615_5020) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1615_5020;
      ov := iv(13 downto 0);
      R_idxprom1615_5024_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5025_root_address_inst
    process(array_obj_ref_5025_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_5025_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_5025_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5108_index_1_rename
    process(R_idxprom1658_5107_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1658_5107_resized;
      ov(13 downto 0) := iv;
      R_idxprom1658_5107_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5108_index_1_resize
    process(idxprom1658_5103) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1658_5103;
      ov := iv(13 downto 0);
      R_idxprom1658_5107_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5108_root_address_inst
    process(array_obj_ref_5108_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_5108_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_5108_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5133_index_1_rename
    process(R_idxprom1663_5132_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1663_5132_resized;
      ov(13 downto 0) := iv;
      R_idxprom1663_5132_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5133_index_1_resize
    process(idxprom1663_5128) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1663_5128;
      ov := iv(13 downto 0);
      R_idxprom1663_5132_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5133_root_address_inst
    process(array_obj_ref_5133_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_5133_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_5133_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1076_addr_0
    process(ptr_deref_1076_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1076_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1076_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1076_base_resize
    process(arrayidx_1074) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1074;
      ov := iv(13 downto 0);
      ptr_deref_1076_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1076_gather_scatter
    process(type_cast_1078_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1078_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1076_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1076_root_address_inst
    process(ptr_deref_1076_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1076_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1076_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1160_addr_0
    process(ptr_deref_1160_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1160_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1160_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1160_base_resize
    process(arrayidx131_1157) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx131_1157;
      ov := iv(13 downto 0);
      ptr_deref_1160_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1160_gather_scatter
    process(ptr_deref_1160_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1160_data_0;
      ov(63 downto 0) := iv;
      tmp132_1161 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1160_root_address_inst
    process(ptr_deref_1160_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1160_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1160_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1184_addr_0
    process(ptr_deref_1184_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1184_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1184_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1184_base_resize
    process(arrayidx136_1182) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx136_1182;
      ov := iv(13 downto 0);
      ptr_deref_1184_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1184_gather_scatter
    process(tmp132_1161) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp132_1161;
      ov(63 downto 0) := iv;
      ptr_deref_1184_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1184_root_address_inst
    process(ptr_deref_1184_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1184_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1184_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1364_addr_0
    process(ptr_deref_1364_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1364_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1364_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1364_base_resize
    process(iNsTr_21_1361) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_21_1361;
      ov := iv(6 downto 0);
      ptr_deref_1364_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1364_gather_scatter
    process(ptr_deref_1364_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1364_data_0;
      ov(31 downto 0) := iv;
      tmp213_1365 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1364_root_address_inst
    process(ptr_deref_1364_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1364_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1364_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1376_addr_0
    process(ptr_deref_1376_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1376_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1376_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1376_base_resize
    process(iNsTr_22_1373) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_22_1373;
      ov := iv(6 downto 0);
      ptr_deref_1376_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1376_gather_scatter
    process(ptr_deref_1376_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1376_data_0;
      ov(31 downto 0) := iv;
      tmp217_1377 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1376_root_address_inst
    process(ptr_deref_1376_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1376_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1376_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1633_addr_0
    process(ptr_deref_1633_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1633_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1633_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1633_base_resize
    process(arrayidx299_1631) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx299_1631;
      ov := iv(13 downto 0);
      ptr_deref_1633_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1633_gather_scatter
    process(type_cast_1635_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1635_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1633_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1633_root_address_inst
    process(ptr_deref_1633_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1633_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1633_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1717_addr_0
    process(ptr_deref_1717_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1717_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1717_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1717_base_resize
    process(arrayidx342_1714) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx342_1714;
      ov := iv(13 downto 0);
      ptr_deref_1717_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1717_gather_scatter
    process(ptr_deref_1717_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1717_data_0;
      ov(63 downto 0) := iv;
      tmp343_1718 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1717_root_address_inst
    process(ptr_deref_1717_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1717_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1717_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1741_addr_0
    process(ptr_deref_1741_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1741_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1741_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1741_base_resize
    process(arrayidx347_1739) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx347_1739;
      ov := iv(13 downto 0);
      ptr_deref_1741_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1741_gather_scatter
    process(tmp343_1718) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp343_1718;
      ov(63 downto 0) := iv;
      ptr_deref_1741_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1741_root_address_inst
    process(ptr_deref_1741_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1741_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1741_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1914_addr_0
    process(ptr_deref_1914_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1914_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1914_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1914_base_resize
    process(iNsTr_37_1911) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_37_1911;
      ov := iv(6 downto 0);
      ptr_deref_1914_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1914_gather_scatter
    process(ptr_deref_1914_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1914_data_0;
      ov(31 downto 0) := iv;
      tmp429_1915 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1914_root_address_inst
    process(ptr_deref_1914_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1914_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1914_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1926_addr_0
    process(ptr_deref_1926_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1926_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1926_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1926_base_resize
    process(iNsTr_38_1923) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_38_1923;
      ov := iv(6 downto 0);
      ptr_deref_1926_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1926_gather_scatter
    process(ptr_deref_1926_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1926_data_0;
      ov(31 downto 0) := iv;
      tmp433_1927 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1926_root_address_inst
    process(ptr_deref_1926_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1926_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1926_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2189_addr_0
    process(ptr_deref_2189_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2189_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2189_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2189_base_resize
    process(arrayidx516_2187) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx516_2187;
      ov := iv(13 downto 0);
      ptr_deref_2189_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2189_gather_scatter
    process(type_cast_2191_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2191_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_2189_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2189_root_address_inst
    process(ptr_deref_2189_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2189_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2189_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2273_addr_0
    process(ptr_deref_2273_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2273_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2273_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2273_base_resize
    process(arrayidx559_2270) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx559_2270;
      ov := iv(13 downto 0);
      ptr_deref_2273_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2273_gather_scatter
    process(ptr_deref_2273_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2273_data_0;
      ov(63 downto 0) := iv;
      tmp560_2274 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2273_root_address_inst
    process(ptr_deref_2273_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2273_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2273_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2297_addr_0
    process(ptr_deref_2297_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2297_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2297_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2297_base_resize
    process(arrayidx564_2295) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx564_2295;
      ov := iv(13 downto 0);
      ptr_deref_2297_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2297_gather_scatter
    process(tmp560_2274) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp560_2274;
      ov(63 downto 0) := iv;
      ptr_deref_2297_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2297_root_address_inst
    process(ptr_deref_2297_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2297_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2297_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2491_addr_0
    process(ptr_deref_2491_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2491_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2491_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2491_base_resize
    process(iNsTr_53_2488) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_53_2488;
      ov := iv(6 downto 0);
      ptr_deref_2491_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2491_gather_scatter
    process(ptr_deref_2491_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2491_data_0;
      ov(31 downto 0) := iv;
      tmp651_2492 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2491_root_address_inst
    process(ptr_deref_2491_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2491_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2491_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2503_addr_0
    process(ptr_deref_2503_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2503_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2503_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2503_base_resize
    process(iNsTr_54_2500) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_54_2500;
      ov := iv(6 downto 0);
      ptr_deref_2503_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2503_gather_scatter
    process(ptr_deref_2503_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2503_data_0;
      ov(31 downto 0) := iv;
      tmp655_2504 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2503_root_address_inst
    process(ptr_deref_2503_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2503_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2503_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2759_addr_0
    process(ptr_deref_2759_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2759_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2759_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2759_base_resize
    process(arrayidx737_2757) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx737_2757;
      ov := iv(13 downto 0);
      ptr_deref_2759_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2759_gather_scatter
    process(type_cast_2761_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2761_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_2759_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2759_root_address_inst
    process(ptr_deref_2759_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2759_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2759_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2843_addr_0
    process(ptr_deref_2843_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2843_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2843_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2843_base_resize
    process(arrayidx780_2840) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx780_2840;
      ov := iv(13 downto 0);
      ptr_deref_2843_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2843_gather_scatter
    process(ptr_deref_2843_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2843_data_0;
      ov(63 downto 0) := iv;
      tmp781_2844 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2843_root_address_inst
    process(ptr_deref_2843_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2843_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2843_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2867_addr_0
    process(ptr_deref_2867_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2867_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2867_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2867_base_resize
    process(arrayidx785_2865) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx785_2865;
      ov := iv(13 downto 0);
      ptr_deref_2867_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2867_gather_scatter
    process(tmp781_2844) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp781_2844;
      ov(63 downto 0) := iv;
      ptr_deref_2867_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2867_root_address_inst
    process(ptr_deref_2867_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2867_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2867_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3040_addr_0
    process(ptr_deref_3040_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3040_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_3040_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3040_base_resize
    process(iNsTr_69_3037) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_69_3037;
      ov := iv(6 downto 0);
      ptr_deref_3040_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3040_gather_scatter
    process(ptr_deref_3040_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3040_data_0;
      ov(31 downto 0) := iv;
      tmp867_3041 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3040_root_address_inst
    process(ptr_deref_3040_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3040_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_3040_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3052_addr_0
    process(ptr_deref_3052_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3052_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_3052_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3052_base_resize
    process(iNsTr_70_3049) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_70_3049;
      ov := iv(6 downto 0);
      ptr_deref_3052_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3052_gather_scatter
    process(ptr_deref_3052_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3052_data_0;
      ov(31 downto 0) := iv;
      tmp871_3053 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3052_root_address_inst
    process(ptr_deref_3052_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3052_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_3052_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3321_addr_0
    process(ptr_deref_3321_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3321_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3321_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3321_base_resize
    process(arrayidx955_3319) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx955_3319;
      ov := iv(13 downto 0);
      ptr_deref_3321_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3321_gather_scatter
    process(type_cast_3323_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3323_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_3321_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3321_root_address_inst
    process(ptr_deref_3321_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3321_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3321_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3405_addr_0
    process(ptr_deref_3405_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3405_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3405_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3405_base_resize
    process(arrayidx998_3402) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx998_3402;
      ov := iv(13 downto 0);
      ptr_deref_3405_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3405_gather_scatter
    process(ptr_deref_3405_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3405_data_0;
      ov(63 downto 0) := iv;
      tmp999_3406 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3405_root_address_inst
    process(ptr_deref_3405_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3405_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3405_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3429_addr_0
    process(ptr_deref_3429_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3429_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3429_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3429_base_resize
    process(arrayidx1003_3427) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1003_3427;
      ov := iv(13 downto 0);
      ptr_deref_3429_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3429_gather_scatter
    process(tmp999_3406) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp999_3406;
      ov(63 downto 0) := iv;
      ptr_deref_3429_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3429_root_address_inst
    process(ptr_deref_3429_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3429_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3429_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3629_addr_0
    process(ptr_deref_3629_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3629_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_3629_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3629_base_resize
    process(iNsTr_85_3626) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_85_3626;
      ov := iv(6 downto 0);
      ptr_deref_3629_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3629_gather_scatter
    process(ptr_deref_3629_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3629_data_0;
      ov(31 downto 0) := iv;
      tmp1091_3630 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3629_root_address_inst
    process(ptr_deref_3629_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3629_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_3629_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3641_addr_0
    process(ptr_deref_3641_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3641_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_3641_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3641_base_resize
    process(iNsTr_86_3638) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_86_3638;
      ov := iv(6 downto 0);
      ptr_deref_3641_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3641_gather_scatter
    process(ptr_deref_3641_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3641_data_0;
      ov(31 downto 0) := iv;
      tmp1095_3642 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3641_root_address_inst
    process(ptr_deref_3641_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3641_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_3641_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3903_addr_0
    process(ptr_deref_3903_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3903_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3903_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3903_base_resize
    process(arrayidx1178_3901) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1178_3901;
      ov := iv(13 downto 0);
      ptr_deref_3903_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3903_gather_scatter
    process(type_cast_3905_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3905_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_3903_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3903_root_address_inst
    process(ptr_deref_3903_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3903_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3903_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3987_addr_0
    process(ptr_deref_3987_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3987_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3987_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3987_base_resize
    process(arrayidx1221_3984) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1221_3984;
      ov := iv(13 downto 0);
      ptr_deref_3987_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3987_gather_scatter
    process(ptr_deref_3987_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3987_data_0;
      ov(63 downto 0) := iv;
      tmp1222_3988 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3987_root_address_inst
    process(ptr_deref_3987_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3987_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3987_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4011_addr_0
    process(ptr_deref_4011_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4011_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4011_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4011_base_resize
    process(arrayidx1226_4009) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1226_4009;
      ov := iv(13 downto 0);
      ptr_deref_4011_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4011_gather_scatter
    process(tmp1222_3988) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp1222_3988;
      ov(63 downto 0) := iv;
      ptr_deref_4011_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4011_root_address_inst
    process(ptr_deref_4011_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4011_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4011_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4196_addr_0
    process(ptr_deref_4196_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4196_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_4196_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4196_base_resize
    process(iNsTr_101_4193) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_101_4193;
      ov := iv(6 downto 0);
      ptr_deref_4196_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4196_gather_scatter
    process(ptr_deref_4196_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4196_data_0;
      ov(31 downto 0) := iv;
      tmp1310_4197 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4196_root_address_inst
    process(ptr_deref_4196_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4196_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_4196_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4208_addr_0
    process(ptr_deref_4208_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4208_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_4208_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4208_base_resize
    process(iNsTr_102_4205) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_102_4205;
      ov := iv(6 downto 0);
      ptr_deref_4208_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4208_gather_scatter
    process(ptr_deref_4208_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4208_data_0;
      ov(31 downto 0) := iv;
      tmp1314_4209 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4208_root_address_inst
    process(ptr_deref_4208_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4208_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_4208_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4465_addr_0
    process(ptr_deref_4465_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4465_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4465_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4465_base_resize
    process(arrayidx1396_4463) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1396_4463;
      ov := iv(13 downto 0);
      ptr_deref_4465_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4465_gather_scatter
    process(type_cast_4467_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_4467_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_4465_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4465_root_address_inst
    process(ptr_deref_4465_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4465_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4465_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4549_addr_0
    process(ptr_deref_4549_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4549_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4549_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4549_base_resize
    process(arrayidx1439_4546) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1439_4546;
      ov := iv(13 downto 0);
      ptr_deref_4549_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4549_gather_scatter
    process(ptr_deref_4549_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4549_data_0;
      ov(63 downto 0) := iv;
      tmp1440_4550 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4549_root_address_inst
    process(ptr_deref_4549_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4549_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4549_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4573_addr_0
    process(ptr_deref_4573_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4573_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4573_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4573_base_resize
    process(arrayidx1444_4571) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1444_4571;
      ov := iv(13 downto 0);
      ptr_deref_4573_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4573_gather_scatter
    process(tmp1440_4550) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp1440_4550;
      ov(63 downto 0) := iv;
      ptr_deref_4573_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4573_root_address_inst
    process(ptr_deref_4573_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4573_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4573_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4767_addr_0
    process(ptr_deref_4767_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4767_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_4767_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4767_base_resize
    process(iNsTr_117_4764) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_117_4764;
      ov := iv(6 downto 0);
      ptr_deref_4767_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4767_gather_scatter
    process(ptr_deref_4767_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4767_data_0;
      ov(31 downto 0) := iv;
      tmp1531_4768 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4767_root_address_inst
    process(ptr_deref_4767_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4767_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_4767_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4779_addr_0
    process(ptr_deref_4779_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4779_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_4779_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4779_base_resize
    process(iNsTr_118_4776) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_118_4776;
      ov := iv(6 downto 0);
      ptr_deref_4779_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4779_gather_scatter
    process(ptr_deref_4779_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4779_data_0;
      ov(31 downto 0) := iv;
      tmp1535_4780 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4779_root_address_inst
    process(ptr_deref_4779_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4779_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_4779_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5029_addr_0
    process(ptr_deref_5029_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5029_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_5029_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5029_base_resize
    process(arrayidx1616_5027) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1616_5027;
      ov := iv(13 downto 0);
      ptr_deref_5029_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5029_gather_scatter
    process(type_cast_5031_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_5031_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_5029_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5029_root_address_inst
    process(ptr_deref_5029_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5029_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_5029_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5113_addr_0
    process(ptr_deref_5113_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5113_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_5113_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5113_base_resize
    process(arrayidx1659_5110) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1659_5110;
      ov := iv(13 downto 0);
      ptr_deref_5113_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5113_gather_scatter
    process(ptr_deref_5113_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5113_data_0;
      ov(63 downto 0) := iv;
      tmp1660_5114 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5113_root_address_inst
    process(ptr_deref_5113_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5113_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_5113_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5137_addr_0
    process(ptr_deref_5137_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5137_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_5137_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5137_base_resize
    process(arrayidx1664_5135) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1664_5135;
      ov := iv(13 downto 0);
      ptr_deref_5137_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5137_gather_scatter
    process(tmp1660_5114) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp1660_5114;
      ov(63 downto 0) := iv;
      ptr_deref_5137_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5137_root_address_inst
    process(ptr_deref_5137_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5137_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_5137_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_727_addr_0
    process(ptr_deref_727_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_727_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_727_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_727_base_resize
    process(iNsTr_0_724) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_724;
      ov := iv(6 downto 0);
      ptr_deref_727_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_727_gather_scatter
    process(ptr_deref_727_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_727_data_0;
      ov(31 downto 0) := iv;
      tmp_728 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_727_root_address_inst
    process(ptr_deref_727_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_727_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_727_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_746_addr_0
    process(ptr_deref_746_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_746_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_746_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_746_base_resize
    process(iNsTr_2_743) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_743;
      ov := iv(6 downto 0);
      ptr_deref_746_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_746_gather_scatter
    process(ptr_deref_746_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_746_data_0;
      ov(31 downto 0) := iv;
      tmp1_747 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_746_root_address_inst
    process(ptr_deref_746_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_746_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_746_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_765_addr_0
    process(ptr_deref_765_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_765_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_765_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_765_base_resize
    process(iNsTr_4_762) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_762;
      ov := iv(6 downto 0);
      ptr_deref_765_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_765_gather_scatter
    process(ptr_deref_765_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_765_data_0;
      ov(31 downto 0) := iv;
      tmp3_766 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_765_root_address_inst
    process(ptr_deref_765_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_765_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_765_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_794_addr_0
    process(ptr_deref_794_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_794_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_794_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_794_base_resize
    process(iNsTr_7_791) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_791;
      ov := iv(6 downto 0);
      ptr_deref_794_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_794_gather_scatter
    process(ptr_deref_794_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_794_data_0;
      ov(31 downto 0) := iv;
      tmp21_795 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_794_root_address_inst
    process(ptr_deref_794_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_794_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_794_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_806_addr_0
    process(ptr_deref_806_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_806_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_806_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_806_base_resize
    process(iNsTr_8_803) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_803;
      ov := iv(6 downto 0);
      ptr_deref_806_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_806_gather_scatter
    process(ptr_deref_806_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_806_data_0;
      ov(31 downto 0) := iv;
      tmp24_807 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_806_root_address_inst
    process(ptr_deref_806_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_806_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_806_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_1016_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp74_1015;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1016_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1016_branch_req_0,
          ack0 => if_stmt_1016_branch_ack_0,
          ack1 => if_stmt_1016_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1207_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp143_1206;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1207_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1207_branch_req_0,
          ack0 => if_stmt_1207_branch_ack_0,
          ack1 => if_stmt_1207_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1300_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp176_1299;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1300_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1300_branch_req_0,
          ack0 => if_stmt_1300_branch_ack_0,
          ack1 => if_stmt_1300_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1497_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp249_1496;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1497_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1497_branch_req_0,
          ack0 => if_stmt_1497_branch_ack_0,
          ack1 => if_stmt_1497_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1529_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp260_1528;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1529_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1529_branch_req_0,
          ack0 => if_stmt_1529_branch_ack_0,
          ack1 => if_stmt_1529_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1548_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp267_1547;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1548_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1548_branch_req_0,
          ack0 => if_stmt_1548_branch_ack_0,
          ack1 => if_stmt_1548_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1574_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp277_1573;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1574_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1574_branch_req_0,
          ack0 => if_stmt_1574_branch_ack_0,
          ack1 => if_stmt_1574_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1764_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp356_1763;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1764_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1764_branch_req_0,
          ack0 => if_stmt_1764_branch_ack_0,
          ack1 => if_stmt_1764_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1850_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp390_1849;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1850_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1850_branch_req_0,
          ack0 => if_stmt_1850_branch_ack_0,
          ack1 => if_stmt_1850_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2047_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp465_2046;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2047_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2047_branch_req_0,
          ack0 => if_stmt_2047_branch_ack_0,
          ack1 => if_stmt_2047_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2079_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp476_2078;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2079_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2079_branch_req_0,
          ack0 => if_stmt_2079_branch_ack_0,
          ack1 => if_stmt_2079_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2098_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp483_2097;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2098_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2098_branch_req_0,
          ack0 => if_stmt_2098_branch_ack_0,
          ack1 => if_stmt_2098_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2130_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp494_2129;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2130_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2130_branch_req_0,
          ack0 => if_stmt_2130_branch_ack_0,
          ack1 => if_stmt_2130_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2320_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp573_2319;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2320_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2320_branch_req_0,
          ack0 => if_stmt_2320_branch_ack_0,
          ack1 => if_stmt_2320_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2413_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp608_2412;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2413_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2413_branch_req_0,
          ack0 => if_stmt_2413_branch_ack_0,
          ack1 => if_stmt_2413_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2623_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp687_2622;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2623_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2623_branch_req_0,
          ack0 => if_stmt_2623_branch_ack_0,
          ack1 => if_stmt_2623_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2655_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp698_2654;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2655_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2655_branch_req_0,
          ack0 => if_stmt_2655_branch_ack_0,
          ack1 => if_stmt_2655_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2674_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp705_2673;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2674_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2674_branch_req_0,
          ack0 => if_stmt_2674_branch_ack_0,
          ack1 => if_stmt_2674_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2700_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp715_2699;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2700_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2700_branch_req_0,
          ack0 => if_stmt_2700_branch_ack_0,
          ack1 => if_stmt_2700_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2890_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp794_2889;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2890_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2890_branch_req_0,
          ack0 => if_stmt_2890_branch_ack_0,
          ack1 => if_stmt_2890_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2976_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp828_2975;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2976_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2976_branch_req_0,
          ack0 => if_stmt_2976_branch_ack_0,
          ack1 => if_stmt_2976_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3173_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp903_3172;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3173_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3173_branch_req_0,
          ack0 => if_stmt_3173_branch_ack_0,
          ack1 => if_stmt_3173_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3211_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp915_3210;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3211_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3211_branch_req_0,
          ack0 => if_stmt_3211_branch_ack_0,
          ack1 => if_stmt_3211_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3230_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp922_3229;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3230_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3230_branch_req_0,
          ack0 => if_stmt_3230_branch_ack_0,
          ack1 => if_stmt_3230_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3262_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp933_3261;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3262_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3262_branch_req_0,
          ack0 => if_stmt_3262_branch_ack_0,
          ack1 => if_stmt_3262_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3452_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1012_3451;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3452_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3452_branch_req_0,
          ack0 => if_stmt_3452_branch_ack_0,
          ack1 => if_stmt_3452_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3551_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1048_3550;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3551_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3551_branch_req_0,
          ack0 => if_stmt_3551_branch_ack_0,
          ack1 => if_stmt_3551_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3761_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1127_3760;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3761_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3761_branch_req_0,
          ack0 => if_stmt_3761_branch_ack_0,
          ack1 => if_stmt_3761_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3799_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1139_3798;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3799_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3799_branch_req_0,
          ack0 => if_stmt_3799_branch_ack_0,
          ack1 => if_stmt_3799_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3818_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1146_3817;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3818_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3818_branch_req_0,
          ack0 => if_stmt_3818_branch_ack_0,
          ack1 => if_stmt_3818_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3844_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1156_3843;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3844_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3844_branch_req_0,
          ack0 => if_stmt_3844_branch_ack_0,
          ack1 => if_stmt_3844_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4034_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1235_4033;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4034_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4034_branch_req_0,
          ack0 => if_stmt_4034_branch_ack_0,
          ack1 => if_stmt_4034_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4126_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1270_4125;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4126_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4126_branch_req_0,
          ack0 => if_stmt_4126_branch_ack_0,
          ack1 => if_stmt_4126_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4329_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1346_4328;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4329_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4329_branch_req_0,
          ack0 => if_stmt_4329_branch_ack_0,
          ack1 => if_stmt_4329_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4355_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1356_4354;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4355_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4355_branch_req_0,
          ack0 => if_stmt_4355_branch_ack_0,
          ack1 => if_stmt_4355_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4374_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1363_4373;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4374_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4374_branch_req_0,
          ack0 => if_stmt_4374_branch_ack_0,
          ack1 => if_stmt_4374_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4406_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1374_4405;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4406_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4406_branch_req_0,
          ack0 => if_stmt_4406_branch_ack_0,
          ack1 => if_stmt_4406_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4596_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1453_4595;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4596_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4596_branch_req_0,
          ack0 => if_stmt_4596_branch_ack_0,
          ack1 => if_stmt_4596_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4683_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1487_4682;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4683_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4683_branch_req_0,
          ack0 => if_stmt_4683_branch_ack_0,
          ack1 => if_stmt_4683_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4899_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1567_4898;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4899_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4899_branch_req_0,
          ack0 => if_stmt_4899_branch_ack_0,
          ack1 => if_stmt_4899_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4925_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1577_4924;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4925_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4925_branch_req_0,
          ack0 => if_stmt_4925_branch_ack_0,
          ack1 => if_stmt_4925_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4944_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1584_4943;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4944_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4944_branch_req_0,
          ack0 => if_stmt_4944_branch_ack_0,
          ack1 => if_stmt_4944_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4970_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1594_4969;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4970_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4970_branch_req_0,
          ack0 => if_stmt_4970_branch_ack_0,
          ack1 => if_stmt_4970_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_5160_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1673_5159;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_5160_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_5160_branch_req_0,
          ack0 => if_stmt_5160_branch_ack_0,
          ack1 => if_stmt_5160_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_5240_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1706_5239;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_5240_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_5240_branch_req_0,
          ack0 => if_stmt_5240_branch_ack_0,
          ack1 => if_stmt_5240_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_933_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_932;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_933_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_933_branch_req_0,
          ack0 => if_stmt_933_branch_ack_0,
          ack1 => if_stmt_933_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_965_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp56_964;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_965_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_965_branch_req_0,
          ack0 => if_stmt_965_branch_ack_0,
          ack1 => if_stmt_965_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_984_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp63_983;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_984_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_984_branch_req_0,
          ack0 => if_stmt_984_branch_ack_0,
          ack1 => if_stmt_984_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1218_inst
    process(kx_x1_913) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_913, type_cast_1217_wire_constant, tmp_var);
      add148_1219 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1226_inst
    process(jx_x1_899) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_899, type_cast_1225_wire_constant, tmp_var);
      inc_1227 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1263_inst
    process(inc165_1259, ix_x2_906) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc165_1259, ix_x2_906, tmp_var);
      inc165x_xix_x2_1264 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1775_inst
    process(k186x_x1_1477) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k186x_x1_1477, type_cast_1774_wire_constant, tmp_var);
      add361_1776 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1783_inst
    process(j240x_x1_1464) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j240x_x1_1464, type_cast_1782_wire_constant, tmp_var);
      inc365_1784 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1814_inst
    process(inc379_1810, i194x_x2_1470) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc379_1810, i194x_x2_1470, tmp_var);
      inc379x_xi194x_x2_1815 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2331_inst
    process(k402x_x1_2014) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k402x_x1_2014, type_cast_2330_wire_constant, tmp_var);
      add578_2332 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2339_inst
    process(j456x_x1_2027) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j456x_x1_2027, type_cast_2338_wire_constant, tmp_var);
      inc582_2340 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2376_inst
    process(inc597_2372, i406x_x2_2021) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc597_2372, i406x_x2_2021, tmp_var);
      inc597x_xi406x_x2_2377 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2901_inst
    process(k620x_x1_2591) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k620x_x1_2591, type_cast_2900_wire_constant, tmp_var);
      add799_2902 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2909_inst
    process(j678x_x1_2604) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j678x_x1_2604, type_cast_2908_wire_constant, tmp_var);
      inc803_2910 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2940_inst
    process(inc817_2936, i628x_x2_2598) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc817_2936, i628x_x2_2598, tmp_var);
      inc817x_xi628x_x2_2941 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3463_inst
    process(k840x_x1_3140) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k840x_x1_3140, type_cast_3462_wire_constant, tmp_var);
      add1017_3464 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3471_inst
    process(j894x_x1_3153) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j894x_x1_3153, type_cast_3470_wire_constant, tmp_var);
      inc1021_3472 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3508_inst
    process(inc1036_3504, i844x_x2_3147) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1036_3504, i844x_x2_3147, tmp_var);
      inc1036x_xi844x_x2_3509 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4045_inst
    process(k1060x_x1_3729) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k1060x_x1_3729, type_cast_4044_wire_constant, tmp_var);
      add1240_4046 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4053_inst
    process(j1118x_x1_3742) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j1118x_x1_3742, type_cast_4052_wire_constant, tmp_var);
      inc1244_4054 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4084_inst
    process(inc1258_4080, i1068x_x2_3736) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1258_4080, i1068x_x2_3736, tmp_var);
      inc1258x_xi1068x_x2_4085 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4607_inst
    process(k1282x_x1_4296) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k1282x_x1_4296, type_cast_4606_wire_constant, tmp_var);
      add1458_4608 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4615_inst
    process(j1337x_x1_4309) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j1337x_x1_4309, type_cast_4614_wire_constant, tmp_var);
      inc1462_4616 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4652_inst
    process(inc1477_4648, i1286x_x2_4303) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1477_4648, i1286x_x2_4303, tmp_var);
      inc1477x_xi1286x_x2_4653 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_5171_inst
    process(k1499x_x1_4867) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k1499x_x1_4867, type_cast_5170_wire_constant, tmp_var);
      add1678_5172 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_5179_inst
    process(j1558x_x1_4880) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j1558x_x1_4880, type_cast_5178_wire_constant, tmp_var);
      inc1682_5180 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_5210_inst
    process(inc1696_5206, i1507x_x2_4874) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1696_5206, i1507x_x2_4874, tmp_var);
      inc1696x_xi1507x_x2_5211 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1007_inst
    process(div70_1003, conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div70_1003, conv48_855, tmp_var);
      add73_1008 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1046_inst
    process(mul89_1042, mul83_1037) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul89_1042, mul83_1037, tmp_var);
      add84_1047 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1051_inst
    process(add84_1047, conv78_1027) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add84_1047, conv78_1027, tmp_var);
      add90_1052 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1110_inst
    process(conv94_1086, mul101_1096) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv94_1086, mul101_1096, tmp_var);
      add102_1111 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1115_inst
    process(add102_1111, mul110_1106) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add102_1111, mul110_1106, tmp_var);
      add111_1116 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1130_inst
    process(mul126_1126, mul120_1121) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul126_1126, mul120_1121, tmp_var);
      add121_1131 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1135_inst
    process(add121_1131, conv94_1086) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add121_1131, conv94_1086, tmp_var);
      add127_1136 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1198_inst
    process(conv139_1193) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv139_1193, type_cast_1197_wire_constant, tmp_var);
      add140_1199 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1249_inst
    process(div156_1245, shl_876) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div156_1245, shl_876, tmp_var);
      add159_1250 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1293_inst
    process(div171_1289, shl_876) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div171_1289, shl_876, tmp_var);
      add175_1294 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1520_inst
    process(div256_1516, conv248_1420) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div256_1516, conv248_1420, tmp_var);
      add259_1521 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1565_inst
    process(conv273_1561, conv248_1420) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv273_1561, conv248_1420, tmp_var);
      add276_1566 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1604_inst
    process(mul294_1600, mul288_1595) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul294_1600, mul288_1595, tmp_var);
      add289_1605 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1609_inst
    process(add289_1605, conv283_1585) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add289_1605, conv283_1585, tmp_var);
      add295_1610 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1667_inst
    process(conv304_1643, mul312_1653) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv304_1643, mul312_1653, tmp_var);
      add313_1668 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1672_inst
    process(add313_1668, mul321_1663) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add313_1668, mul321_1663, tmp_var);
      add322_1673 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1687_inst
    process(mul337_1683, mul331_1678) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul337_1683, mul331_1678, tmp_var);
      add332_1688 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1692_inst
    process(add332_1688, conv304_1643) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add332_1688, conv304_1643, tmp_var);
      add338_1693 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1755_inst
    process(conv352_1750) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv352_1750, type_cast_1754_wire_constant, tmp_var);
      add353_1756 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1800_inst
    process(conv369_1796, shl372_1441) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv369_1796, shl372_1441, tmp_var);
      add373_1801 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1843_inst
    process(div385_1839, shl372_1441) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div385_1839, shl372_1441, tmp_var);
      add389_1844 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2070_inst
    process(div472_2066, conv464_1970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div472_2066, conv464_1970, tmp_var);
      add475_2071 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2121_inst
    process(div490_2117, conv464_1970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div490_2117, conv464_1970, tmp_var);
      add493_2122 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2160_inst
    process(mul511_2156, conv500_2141) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul511_2156, conv500_2141, tmp_var);
      add506_2161 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2165_inst
    process(add506_2161, mul505_2151) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add506_2161, mul505_2151, tmp_var);
      add512_2166 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2223_inst
    process(mul538_2219, conv521_2199) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul538_2219, conv521_2199, tmp_var);
      add530_2224 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2228_inst
    process(add530_2224, mul529_2209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add530_2224, mul529_2209, tmp_var);
      add539_2229 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2243_inst
    process(mul554_2239, conv521_2199) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul554_2239, conv521_2199, tmp_var);
      add549_2244 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2248_inst
    process(add549_2244, mul548_2234) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add549_2244, mul548_2234, tmp_var);
      add555_2249 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2311_inst
    process(conv569_2306) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv569_2306, type_cast_2310_wire_constant, tmp_var);
      add570_2312 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2362_inst
    process(div587_2358, shl590_1991) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div587_2358, shl590_1991, tmp_var);
      add591_2363 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2406_inst
    process(div603_2402, shl590_1991) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div603_2402, shl590_1991, tmp_var);
      add607_2407 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2646_inst
    process(div694_2642, conv686_2547) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div694_2642, conv686_2547, tmp_var);
      add697_2647 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2691_inst
    process(conv711_2687, conv686_2547) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv711_2687, conv686_2547, tmp_var);
      add714_2692 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2730_inst
    process(mul732_2726, conv721_2711) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul732_2726, conv721_2711, tmp_var);
      add727_2731 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2735_inst
    process(add727_2731, mul726_2721) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add727_2731, mul726_2721, tmp_var);
      add733_2736 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2793_inst
    process(mul759_2789, conv742_2769) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul759_2789, conv742_2769, tmp_var);
      add751_2794 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2798_inst
    process(add751_2794, mul750_2779) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add751_2794, mul750_2779, tmp_var);
      add760_2799 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2813_inst
    process(mul775_2809, conv742_2769) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul775_2809, conv742_2769, tmp_var);
      add770_2814 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2818_inst
    process(add770_2814, mul769_2804) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add770_2814, mul769_2804, tmp_var);
      add776_2819 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2881_inst
    process(conv790_2876) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv790_2876, type_cast_2880_wire_constant, tmp_var);
      add791_2882 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2926_inst
    process(conv807_2922, shl810_2568) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv807_2922, shl810_2568, tmp_var);
      add811_2927 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2969_inst
    process(div823_2965, shl810_2568) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div823_2965, shl810_2568, tmp_var);
      add827_2970 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3202_inst
    process(div911_3198, conv902_3096) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div911_3198, conv902_3096, tmp_var);
      add914_3203 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3253_inst
    process(div929_3249, conv902_3096) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div929_3249, conv902_3096, tmp_var);
      add932_3254 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3292_inst
    process(mul950_3288, conv939_3273) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul950_3288, conv939_3273, tmp_var);
      add945_3293 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3297_inst
    process(add945_3293, mul944_3283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add945_3293, mul944_3283, tmp_var);
      add951_3298 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3355_inst
    process(mul977_3351, conv960_3331) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul977_3351, conv960_3331, tmp_var);
      add969_3356 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3360_inst
    process(add969_3356, mul968_3341) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add969_3356, mul968_3341, tmp_var);
      add978_3361 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3375_inst
    process(mul993_3371, conv960_3331) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul993_3371, conv960_3331, tmp_var);
      add988_3376 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3380_inst
    process(add988_3376, mul987_3366) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add988_3376, mul987_3366, tmp_var);
      add994_3381 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3443_inst
    process(conv1008_3438) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1008_3438, type_cast_3442_wire_constant, tmp_var);
      add1009_3444 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3494_inst
    process(div1026_3490, shl1029_3117) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1026_3490, shl1029_3117, tmp_var);
      add1030_3495 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3544_inst
    process(div1043_3540, shl1029_3117) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1043_3540, shl1029_3117, tmp_var);
      add1047_3545 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3790_inst
    process(div1135_3786, conv1126_3685) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1135_3786, conv1126_3685, tmp_var);
      add1138_3791 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3835_inst
    process(conv1152_3831, conv1126_3685) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1152_3831, conv1126_3685, tmp_var);
      add1155_3836 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3874_inst
    process(mul1173_3870, conv1162_3855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1173_3870, conv1162_3855, tmp_var);
      add1168_3875 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3879_inst
    process(add1168_3875, mul1167_3865) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1168_3875, mul1167_3865, tmp_var);
      add1174_3880 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3937_inst
    process(mul1200_3933, conv1183_3913) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1200_3933, conv1183_3913, tmp_var);
      add1192_3938 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3942_inst
    process(add1192_3938, mul1191_3923) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1192_3938, mul1191_3923, tmp_var);
      add1201_3943 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3957_inst
    process(mul1216_3953, conv1183_3913) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1216_3953, conv1183_3913, tmp_var);
      add1211_3958 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3962_inst
    process(add1211_3958, mul1210_3948) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1211_3958, mul1210_3948, tmp_var);
      add1217_3963 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4025_inst
    process(conv1231_4020) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1231_4020, type_cast_4024_wire_constant, tmp_var);
      add1232_4026 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4070_inst
    process(conv1248_4066, shl1251_3706) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1248_4066, shl1251_3706, tmp_var);
      add1252_4071 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4119_inst
    process(div1265_4115, shl1251_3706) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1265_4115, shl1251_3706, tmp_var);
      add1269_4120 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4346_inst
    process(conv1352_4342, conv1345_4252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1352_4342, conv1345_4252, tmp_var);
      add1355_4347 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4397_inst
    process(div1370_4393, conv1345_4252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1370_4393, conv1345_4252, tmp_var);
      add1373_4398 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4436_inst
    process(mul1391_4432, conv1380_4417) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1391_4432, conv1380_4417, tmp_var);
      add1386_4437 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4441_inst
    process(add1386_4437, mul1385_4427) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1386_4437, mul1385_4427, tmp_var);
      add1392_4442 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4499_inst
    process(mul1418_4495, conv1401_4475) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1418_4495, conv1401_4475, tmp_var);
      add1410_4500 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4504_inst
    process(add1410_4500, mul1409_4485) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1410_4500, mul1409_4485, tmp_var);
      add1419_4505 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4519_inst
    process(mul1434_4515, conv1401_4475) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1434_4515, conv1401_4475, tmp_var);
      add1429_4520 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4524_inst
    process(add1429_4520, mul1428_4510) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1429_4520, mul1428_4510, tmp_var);
      add1435_4525 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4587_inst
    process(conv1449_4582) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1449_4582, type_cast_4586_wire_constant, tmp_var);
      add1450_4588 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4638_inst
    process(div1467_4634, shl1470_4273) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1467_4634, shl1470_4273, tmp_var);
      add1471_4639 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4676_inst
    process(conv1482_4672, shl1470_4273) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1482_4672, shl1470_4273, tmp_var);
      add1486_4677 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4916_inst
    process(conv1573_4912, conv1566_4823) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1573_4912, conv1566_4823, tmp_var);
      add1576_4917 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4961_inst
    process(conv1590_4957, conv1566_4823) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1590_4957, conv1566_4823, tmp_var);
      add1593_4962 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5000_inst
    process(mul1611_4996, conv1600_4981) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1611_4996, conv1600_4981, tmp_var);
      add1606_5001 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5005_inst
    process(add1606_5001, mul1605_4991) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1606_5001, mul1605_4991, tmp_var);
      add1612_5006 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5063_inst
    process(mul1638_5059, conv1621_5039) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1638_5059, conv1621_5039, tmp_var);
      add1630_5064 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5068_inst
    process(add1630_5064, mul1629_5049) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1630_5064, mul1629_5049, tmp_var);
      add1639_5069 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5083_inst
    process(mul1654_5079, conv1621_5039) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1654_5079, conv1621_5039, tmp_var);
      add1649_5084 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5088_inst
    process(add1649_5084, mul1648_5074) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1649_5084, mul1648_5074, tmp_var);
      add1655_5089 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5151_inst
    process(conv1669_5146) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1669_5146, type_cast_5150_wire_constant, tmp_var);
      add1670_5152 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5196_inst
    process(conv1686_5192, shl1689_4844) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1686_5192, shl1689_4844, tmp_var);
      add1690_5197 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5233_inst
    process(conv1701_5229, shl1689_4844) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1701_5229, shl1689_4844, tmp_var);
      add1705_5234 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_956_inst
    process(div_952, conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div_952, conv48_855, tmp_var);
      add_957 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1059_inst
    process(type_cast_1055_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1055_wire, type_cast_1058_wire_constant, tmp_var);
      ASHR_i32_i32_1059_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1143_inst
    process(type_cast_1139_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1139_wire, type_cast_1142_wire_constant, tmp_var);
      ASHR_i32_i32_1143_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1168_inst
    process(type_cast_1164_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1164_wire, type_cast_1167_wire_constant, tmp_var);
      ASHR_i32_i32_1168_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1394_inst
    process(type_cast_1390_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1390_wire, type_cast_1393_wire_constant, tmp_var);
      ASHR_i32_i32_1394_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1409_inst
    process(type_cast_1405_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1405_wire, type_cast_1408_wire_constant, tmp_var);
      ASHR_i32_i32_1409_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1433_inst
    process(type_cast_1429_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1429_wire, type_cast_1432_wire_constant, tmp_var);
      ASHR_i32_i32_1433_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1459_inst
    process(type_cast_1455_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1455_wire, type_cast_1458_wire_constant, tmp_var);
      ASHR_i32_i32_1459_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1617_inst
    process(type_cast_1613_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1613_wire, type_cast_1616_wire_constant, tmp_var);
      ASHR_i32_i32_1617_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1700_inst
    process(type_cast_1696_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1696_wire, type_cast_1699_wire_constant, tmp_var);
      ASHR_i32_i32_1700_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1725_inst
    process(type_cast_1721_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1721_wire, type_cast_1724_wire_constant, tmp_var);
      ASHR_i32_i32_1725_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1944_inst
    process(type_cast_1940_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1940_wire, type_cast_1943_wire_constant, tmp_var);
      ASHR_i32_i32_1944_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1959_inst
    process(type_cast_1955_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1955_wire, type_cast_1958_wire_constant, tmp_var);
      ASHR_i32_i32_1959_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1983_inst
    process(type_cast_1979_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1979_wire, type_cast_1982_wire_constant, tmp_var);
      ASHR_i32_i32_1983_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2009_inst
    process(type_cast_2005_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2005_wire, type_cast_2008_wire_constant, tmp_var);
      ASHR_i32_i32_2009_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2173_inst
    process(type_cast_2169_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2169_wire, type_cast_2172_wire_constant, tmp_var);
      ASHR_i32_i32_2173_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2256_inst
    process(type_cast_2252_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2252_wire, type_cast_2255_wire_constant, tmp_var);
      ASHR_i32_i32_2256_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2281_inst
    process(type_cast_2277_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2277_wire, type_cast_2280_wire_constant, tmp_var);
      ASHR_i32_i32_2281_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2521_inst
    process(type_cast_2517_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2517_wire, type_cast_2520_wire_constant, tmp_var);
      ASHR_i32_i32_2521_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2536_inst
    process(type_cast_2532_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2532_wire, type_cast_2535_wire_constant, tmp_var);
      ASHR_i32_i32_2536_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2560_inst
    process(type_cast_2556_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2556_wire, type_cast_2559_wire_constant, tmp_var);
      ASHR_i32_i32_2560_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2586_inst
    process(type_cast_2582_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2582_wire, type_cast_2585_wire_constant, tmp_var);
      ASHR_i32_i32_2586_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2743_inst
    process(type_cast_2739_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2739_wire, type_cast_2742_wire_constant, tmp_var);
      ASHR_i32_i32_2743_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2826_inst
    process(type_cast_2822_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2822_wire, type_cast_2825_wire_constant, tmp_var);
      ASHR_i32_i32_2826_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2851_inst
    process(type_cast_2847_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2847_wire, type_cast_2850_wire_constant, tmp_var);
      ASHR_i32_i32_2851_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3070_inst
    process(type_cast_3066_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3066_wire, type_cast_3069_wire_constant, tmp_var);
      ASHR_i32_i32_3070_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3085_inst
    process(type_cast_3081_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3081_wire, type_cast_3084_wire_constant, tmp_var);
      ASHR_i32_i32_3085_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3109_inst
    process(type_cast_3105_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3105_wire, type_cast_3108_wire_constant, tmp_var);
      ASHR_i32_i32_3109_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3135_inst
    process(type_cast_3131_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3131_wire, type_cast_3134_wire_constant, tmp_var);
      ASHR_i32_i32_3135_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3305_inst
    process(type_cast_3301_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3301_wire, type_cast_3304_wire_constant, tmp_var);
      ASHR_i32_i32_3305_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3388_inst
    process(type_cast_3384_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3384_wire, type_cast_3387_wire_constant, tmp_var);
      ASHR_i32_i32_3388_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3413_inst
    process(type_cast_3409_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3409_wire, type_cast_3412_wire_constant, tmp_var);
      ASHR_i32_i32_3413_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3659_inst
    process(type_cast_3655_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3655_wire, type_cast_3658_wire_constant, tmp_var);
      ASHR_i32_i32_3659_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3674_inst
    process(type_cast_3670_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3670_wire, type_cast_3673_wire_constant, tmp_var);
      ASHR_i32_i32_3674_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3698_inst
    process(type_cast_3694_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3694_wire, type_cast_3697_wire_constant, tmp_var);
      ASHR_i32_i32_3698_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3724_inst
    process(type_cast_3720_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3720_wire, type_cast_3723_wire_constant, tmp_var);
      ASHR_i32_i32_3724_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3887_inst
    process(type_cast_3883_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3883_wire, type_cast_3886_wire_constant, tmp_var);
      ASHR_i32_i32_3887_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3970_inst
    process(type_cast_3966_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3966_wire, type_cast_3969_wire_constant, tmp_var);
      ASHR_i32_i32_3970_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3995_inst
    process(type_cast_3991_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3991_wire, type_cast_3994_wire_constant, tmp_var);
      ASHR_i32_i32_3995_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4226_inst
    process(type_cast_4222_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4222_wire, type_cast_4225_wire_constant, tmp_var);
      ASHR_i32_i32_4226_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4241_inst
    process(type_cast_4237_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4237_wire, type_cast_4240_wire_constant, tmp_var);
      ASHR_i32_i32_4241_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4265_inst
    process(type_cast_4261_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4261_wire, type_cast_4264_wire_constant, tmp_var);
      ASHR_i32_i32_4265_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4291_inst
    process(type_cast_4287_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4287_wire, type_cast_4290_wire_constant, tmp_var);
      ASHR_i32_i32_4291_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4449_inst
    process(type_cast_4445_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4445_wire, type_cast_4448_wire_constant, tmp_var);
      ASHR_i32_i32_4449_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4532_inst
    process(type_cast_4528_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4528_wire, type_cast_4531_wire_constant, tmp_var);
      ASHR_i32_i32_4532_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4557_inst
    process(type_cast_4553_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4553_wire, type_cast_4556_wire_constant, tmp_var);
      ASHR_i32_i32_4557_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4797_inst
    process(type_cast_4793_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4793_wire, type_cast_4796_wire_constant, tmp_var);
      ASHR_i32_i32_4797_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4812_inst
    process(type_cast_4808_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4808_wire, type_cast_4811_wire_constant, tmp_var);
      ASHR_i32_i32_4812_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4836_inst
    process(type_cast_4832_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4832_wire, type_cast_4835_wire_constant, tmp_var);
      ASHR_i32_i32_4836_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4862_inst
    process(type_cast_4858_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4858_wire, type_cast_4861_wire_constant, tmp_var);
      ASHR_i32_i32_4862_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_5013_inst
    process(type_cast_5009_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_5009_wire, type_cast_5012_wire_constant, tmp_var);
      ASHR_i32_i32_5013_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_5096_inst
    process(type_cast_5092_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_5092_wire, type_cast_5095_wire_constant, tmp_var);
      ASHR_i32_i32_5096_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_5121_inst
    process(type_cast_5117_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_5117_wire, type_cast_5120_wire_constant, tmp_var);
      ASHR_i32_i32_5121_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_829_inst
    process(type_cast_825_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_825_wire, type_cast_828_wire_constant, tmp_var);
      ASHR_i32_i32_829_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_844_inst
    process(type_cast_840_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_840_wire, type_cast_843_wire_constant, tmp_var);
      ASHR_i32_i32_844_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_868_inst
    process(type_cast_864_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_864_wire, type_cast_867_wire_constant, tmp_var);
      ASHR_i32_i32_868_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_894_inst
    process(type_cast_890_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_890_wire, type_cast_893_wire_constant, tmp_var);
      ASHR_i32_i32_894_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1254_inst
    process(conv153_1232, add159_1250) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv153_1232, add159_1250, tmp_var);
      cmp160_1255 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1298_inst
    process(conv168_1276, add175_1294) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv168_1276, add175_1294, tmp_var);
      cmp176_1299 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1805_inst
    process(conv367_1789, add373_1801) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv367_1789, add373_1801, tmp_var);
      cmp374_1806 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1848_inst
    process(conv382_1826, add389_1844) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv382_1826, add389_1844, tmp_var);
      cmp390_1849 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2367_inst
    process(conv584_2345, add591_2363) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv584_2345, add591_2363, tmp_var);
      cmp592_2368 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2411_inst
    process(conv600_2389, add607_2407) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv600_2389, add607_2407, tmp_var);
      cmp608_2412 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2931_inst
    process(conv805_2915, add811_2927) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv805_2915, add811_2927, tmp_var);
      cmp812_2932 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2974_inst
    process(conv820_2952, add827_2970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv820_2952, add827_2970, tmp_var);
      cmp828_2975 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3499_inst
    process(conv1023_3477, add1030_3495) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1023_3477, add1030_3495, tmp_var);
      cmp1031_3500 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3549_inst
    process(conv1039_3521, add1047_3545) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1039_3521, add1047_3545, tmp_var);
      cmp1048_3550 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4075_inst
    process(conv1246_4059, add1252_4071) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1246_4059, add1252_4071, tmp_var);
      cmp1253_4076 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4124_inst
    process(conv1261_4096, add1269_4120) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1261_4096, add1269_4120, tmp_var);
      cmp1270_4125 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4643_inst
    process(conv1464_4621, add1471_4639) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1464_4621, add1471_4639, tmp_var);
      cmp1472_4644 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4681_inst
    process(conv1480_4665, add1486_4677) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1480_4665, add1486_4677, tmp_var);
      cmp1487_4682 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_5201_inst
    process(conv1684_5185, add1690_5197) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1684_5185, add1690_5197, tmp_var);
      cmp1691_5202 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_5238_inst
    process(conv1699_5222, add1705_5234) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1699_5222, add1705_5234, tmp_var);
      cmp1706_5239 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1346_inst
    process(conv190_1341) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv190_1341, type_cast_1345_wire_constant, tmp_var);
      div191_1347 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1896_inst
    process(conv408_1891) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv408_1891, type_cast_1895_wire_constant, tmp_var);
      div409_1897 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2463_inst
    process(conv624_2458) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv624_2458, type_cast_2462_wire_constant, tmp_var);
      div625_2464 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2473_inst
    process(conv630_2468) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv630_2468, type_cast_2472_wire_constant, tmp_var);
      div631_2474 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3022_inst
    process(conv846_3017) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv846_3017, type_cast_3021_wire_constant, tmp_var);
      div847_3023 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3601_inst
    process(conv1064_3596) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1064_3596, type_cast_3600_wire_constant, tmp_var);
      div1065_3602 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3611_inst
    process(conv1070_3606) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1070_3606, type_cast_3610_wire_constant, tmp_var);
      div1071_3612 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_4172_inst
    process(conv1288_4167) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1288_4167, type_cast_4171_wire_constant, tmp_var);
      div1289_4173 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_4733_inst
    process(conv1503_4728) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1503_4728, type_cast_4732_wire_constant, tmp_var);
      div1504_4734 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_4749_inst
    process(mul1510_4744) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1510_4744, type_cast_4748_wire_constant, tmp_var);
      div1511_4750 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1002_inst
    process(conv69_997) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv69_997, type_cast_1001_wire_constant, tmp_var);
      div70_1003 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1244_inst
    process(conv155_1239) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv155_1239, type_cast_1243_wire_constant, tmp_var);
      div156_1245 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1288_inst
    process(conv170_1283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv170_1283, type_cast_1287_wire_constant, tmp_var);
      div171_1289 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1515_inst
    process(conv255_1510) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv255_1510, type_cast_1514_wire_constant, tmp_var);
      div256_1516 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1838_inst
    process(conv384_1833) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv384_1833, type_cast_1837_wire_constant, tmp_var);
      div385_1839 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2065_inst
    process(conv471_2060) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv471_2060, type_cast_2064_wire_constant, tmp_var);
      div472_2066 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2116_inst
    process(conv489_2111) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv489_2111, type_cast_2115_wire_constant, tmp_var);
      div490_2117 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2357_inst
    process(conv586_2352) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv586_2352, type_cast_2356_wire_constant, tmp_var);
      div587_2358 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2401_inst
    process(conv602_2396) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv602_2396, type_cast_2400_wire_constant, tmp_var);
      div603_2402 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2641_inst
    process(conv693_2636) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv693_2636, type_cast_2640_wire_constant, tmp_var);
      div694_2642 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2964_inst
    process(conv822_2959) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv822_2959, type_cast_2963_wire_constant, tmp_var);
      div823_2965 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3197_inst
    process(mul910_3192) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul910_3192, type_cast_3196_wire_constant, tmp_var);
      div911_3198 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3248_inst
    process(conv928_3243) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv928_3243, type_cast_3247_wire_constant, tmp_var);
      div929_3249 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3489_inst
    process(conv1025_3484) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1025_3484, type_cast_3488_wire_constant, tmp_var);
      div1026_3490 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3539_inst
    process(mul1042_3534) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1042_3534, type_cast_3538_wire_constant, tmp_var);
      div1043_3540 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3785_inst
    process(mul1134_3780) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1134_3780, type_cast_3784_wire_constant, tmp_var);
      div1135_3786 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_4114_inst
    process(mul1264_4109) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1264_4109, type_cast_4113_wire_constant, tmp_var);
      div1265_4115 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_4392_inst
    process(conv1369_4387) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1369_4387, type_cast_4391_wire_constant, tmp_var);
      div1370_4393 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_4633_inst
    process(conv1466_4628) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1466_4628, type_cast_4632_wire_constant, tmp_var);
      div1467_4634 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_951_inst
    process(conv53_946) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv53_946, type_cast_950_wire_constant, tmp_var);
      div_952 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_4178_inst
    process(div1289_4173) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(div1289_4173, type_cast_4177_wire_constant, tmp_var);
      mul1290_4179 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_4743_inst
    process(conv1509_4738) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1509_4738, type_cast_4742_wire_constant, tmp_var);
      mul1510_4744 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1036_inst
    process(conv82_1032, conv37_831) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv82_1032, conv37_831, tmp_var);
      mul83_1037 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1041_inst
    process(conv46_925, conv86_870) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv46_925, conv86_870, tmp_var);
      mul89_1042 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1095_inst
    process(sub_1091, conv31_811) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_1091, conv31_811, tmp_var);
      mul101_1096 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1105_inst
    process(sub109_1101, conv104_896) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub109_1101, conv104_896, tmp_var);
      mul110_1106 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1120_inst
    process(conv60_976, conv37_831) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv60_976, conv37_831, tmp_var);
      mul120_1121 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1125_inst
    process(conv46_925, conv86_870) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv46_925, conv86_870, tmp_var);
      mul126_1126 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1415_inst
    process(conv236_1411, conv234_1396) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv236_1411, conv234_1396, tmp_var);
      mul237_1416 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1451_inst
    process(mul229_1447, conv226_1381) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul229_1447, conv226_1381, tmp_var);
      sext1719_1452 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1594_inst
    process(conv287_1590, conv234_1396) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv287_1590, conv234_1396, tmp_var);
      mul288_1595 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1599_inst
    process(conv246_1489, conv291_1435) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv246_1489, conv291_1435, tmp_var);
      mul294_1600 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1652_inst
    process(sub311_1648, conv226_1381) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub311_1648, conv226_1381, tmp_var);
      mul312_1653 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1662_inst
    process(sub320_1658, conv315_1461) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub320_1658, conv315_1461, tmp_var);
      mul321_1663 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1677_inst
    process(conv264_1540, conv234_1396) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv264_1540, conv234_1396, tmp_var);
      mul331_1678 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1682_inst
    process(conv246_1489, conv291_1435) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv246_1489, conv291_1435, tmp_var);
      mul337_1683 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1965_inst
    process(conv452_1961, conv450_1946) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv452_1961, conv450_1946, tmp_var);
      mul453_1966 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2001_inst
    process(mul445_1997, conv369x_xlcssa_1883) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul445_1997, conv369x_xlcssa_1883, tmp_var);
      sext1721_2002 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2150_inst
    process(conv504_2146, conv450_1946) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv504_2146, conv450_1946, tmp_var);
      mul505_2151 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2155_inst
    process(conv462_2039, conv508_1985) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv462_2039, conv508_1985, tmp_var);
      mul511_2156 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2208_inst
    process(sub528_2204, conv442_1931) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub528_2204, conv442_1931, tmp_var);
      mul529_2209 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2218_inst
    process(sub537_2214, conv532_2011) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub537_2214, conv532_2011, tmp_var);
      mul538_2219 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2233_inst
    process(conv480_2090, conv450_1946) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv480_2090, conv450_1946, tmp_var);
      mul548_2234 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2238_inst
    process(conv462_2039, conv508_1985) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv462_2039, conv508_1985, tmp_var);
      mul554_2239 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2542_inst
    process(conv674_2538, conv672_2523) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv674_2538, conv672_2523, tmp_var);
      mul675_2543 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2578_inst
    process(mul667_2574, conv586x_xlcssa_2446) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul667_2574, conv586x_xlcssa_2446, tmp_var);
      sext1723_2579 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2720_inst
    process(conv725_2716, conv672_2523) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv725_2716, conv672_2523, tmp_var);
      mul726_2721 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2725_inst
    process(conv684_2615, conv729_2562) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv684_2615, conv729_2562, tmp_var);
      mul732_2726 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2778_inst
    process(sub749_2774, conv664_2508) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub749_2774, conv664_2508, tmp_var);
      mul750_2779 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2788_inst
    process(sub758_2784, conv753_2588) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub758_2784, conv753_2588, tmp_var);
      mul759_2789 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2803_inst
    process(conv702_2666, conv672_2523) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv702_2666, conv672_2523, tmp_var);
      mul769_2804 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2808_inst
    process(conv684_2615, conv729_2562) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv684_2615, conv729_2562, tmp_var);
      mul775_2809 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3091_inst
    process(conv890_3087, conv888_3072) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv890_3087, conv888_3072, tmp_var);
      mul891_3092 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3127_inst
    process(mul883_3123, conv807x_xlcssa_3009) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul883_3123, conv807x_xlcssa_3009, tmp_var);
      sext1725_3128 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3191_inst
    process(conv909_3186) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv909_3186, type_cast_3190_wire_constant, tmp_var);
      mul910_3192 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3282_inst
    process(conv943_3278, conv888_3072) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv943_3278, conv888_3072, tmp_var);
      mul944_3283 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3287_inst
    process(conv900_3165, conv947_3111) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv900_3165, conv947_3111, tmp_var);
      mul950_3288 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3340_inst
    process(sub967_3336, conv880_3057) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub967_3336, conv880_3057, tmp_var);
      mul968_3341 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3350_inst
    process(sub976_3346, conv971_3137) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub976_3346, conv971_3137, tmp_var);
      mul977_3351 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3365_inst
    process(conv919_3222, conv888_3072) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv919_3222, conv888_3072, tmp_var);
      mul987_3366 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3370_inst
    process(conv900_3165, conv947_3111) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv900_3165, conv947_3111, tmp_var);
      mul993_3371 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3533_inst
    process(conv1041_3528) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1041_3528, type_cast_3532_wire_constant, tmp_var);
      mul1042_3534 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3680_inst
    process(conv1114_3676, conv1112_3661) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1114_3676, conv1112_3661, tmp_var);
      mul1115_3681 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3716_inst
    process(mul1107_3712, conv1025x_xlcssa_3584) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul1107_3712, conv1025x_xlcssa_3584, tmp_var);
      sext1727_3717 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3779_inst
    process(conv1133_3774) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1133_3774, type_cast_3778_wire_constant, tmp_var);
      mul1134_3780 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3864_inst
    process(conv1166_3860, conv1112_3661) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1166_3860, conv1112_3661, tmp_var);
      mul1167_3865 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3869_inst
    process(conv1124_3753, conv1170_3700) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1124_3753, conv1170_3700, tmp_var);
      mul1173_3870 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3922_inst
    process(sub1190_3918, conv1104_3646) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1190_3918, conv1104_3646, tmp_var);
      mul1191_3923 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3932_inst
    process(sub1199_3928, conv1194_3726) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1199_3928, conv1194_3726, tmp_var);
      mul1200_3933 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3947_inst
    process(conv1143_3810, conv1112_3661) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1143_3810, conv1112_3661, tmp_var);
      mul1210_3948 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3952_inst
    process(conv1124_3753, conv1170_3700) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1124_3753, conv1170_3700, tmp_var);
      mul1216_3953 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4108_inst
    process(conv1263_4103) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1263_4103, type_cast_4107_wire_constant, tmp_var);
      mul1264_4109 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4247_inst
    process(conv1333_4243, conv1331_4228) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1333_4243, conv1331_4228, tmp_var);
      mul1334_4248 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4283_inst
    process(mul1326_4279, conv1248x_xlcssa_4159) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul1326_4279, conv1248x_xlcssa_4159, tmp_var);
      sext1729_4284 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4426_inst
    process(conv1384_4422, conv1331_4228) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1384_4422, conv1331_4228, tmp_var);
      mul1385_4427 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4431_inst
    process(conv1343_4321, conv1388_4267) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1343_4321, conv1388_4267, tmp_var);
      mul1391_4432 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4484_inst
    process(sub1408_4480, conv1323_4213) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1408_4480, conv1323_4213, tmp_var);
      mul1409_4485 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4494_inst
    process(sub1417_4490, conv1412_4293) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1417_4490, conv1412_4293, tmp_var);
      mul1418_4495 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4509_inst
    process(conv1360_4366, conv1331_4228) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1360_4366, conv1331_4228, tmp_var);
      mul1428_4510 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4514_inst
    process(conv1343_4321, conv1388_4267) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1343_4321, conv1388_4267, tmp_var);
      mul1434_4515 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4818_inst
    process(conv1554_4814, conv1552_4799) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1554_4814, conv1552_4799, tmp_var);
      mul1555_4819 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4854_inst
    process(mul1547_4850, conv1466x_xlcssa_4716) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul1547_4850, conv1466x_xlcssa_4716, tmp_var);
      sext1731_4855 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4990_inst
    process(conv1604_4986, conv1552_4799) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1604_4986, conv1552_4799, tmp_var);
      mul1605_4991 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4995_inst
    process(conv1564_4891, conv1608_4838) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1564_4891, conv1608_4838, tmp_var);
      mul1611_4996 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_5048_inst
    process(sub1628_5044, conv1544_4784) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1628_5044, conv1544_4784, tmp_var);
      mul1629_5049 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_5058_inst
    process(sub1637_5054, conv1632_4864) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1637_5054, conv1632_4864, tmp_var);
      mul1638_5059 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_5073_inst
    process(conv1581_4936, conv1552_4799) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1581_4936, conv1552_4799, tmp_var);
      mul1648_5074 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_5078_inst
    process(conv1564_4891, conv1608_4838) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1564_4891, conv1608_4838, tmp_var);
      mul1654_5079 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_850_inst
    process(conv39_846, conv37_831) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv39_846, conv37_831, tmp_var);
      mul40_851 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_886_inst
    process(mul_882, conv33_815) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_882, conv33_815, tmp_var);
      sext1717_887 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1386_inst
    process(tmp213_1365) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp213_1365, type_cast_1385_wire_constant, tmp_var);
      sext1766_1387 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1401_inst
    process(tmp217_1377) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp217_1377, type_cast_1400_wire_constant, tmp_var);
      sext1718_1402 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1425_inst
    process(mul237_1416) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul237_1416, type_cast_1424_wire_constant, tmp_var);
      sext1767_1426 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1440_inst
    process(conv248_1420) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv248_1420, type_cast_1439_wire_constant, tmp_var);
      shl372_1441 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1446_inst
    process(conv155x_xlcssa_1329) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv155x_xlcssa_1329, type_cast_1445_wire_constant, tmp_var);
      mul229_1447 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1936_inst
    process(tmp429_1915) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp429_1915, type_cast_1935_wire_constant, tmp_var);
      sext1768_1937 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1951_inst
    process(tmp433_1927) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp433_1927, type_cast_1950_wire_constant, tmp_var);
      sext1720_1952 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1975_inst
    process(mul453_1966) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul453_1966, type_cast_1974_wire_constant, tmp_var);
      sext1769_1976 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1990_inst
    process(conv464_1970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv464_1970, type_cast_1989_wire_constant, tmp_var);
      shl590_1991 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1996_inst
    process(conv442_1931) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv442_1931, type_cast_1995_wire_constant, tmp_var);
      mul445_1997 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2513_inst
    process(tmp651_2492) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp651_2492, type_cast_2512_wire_constant, tmp_var);
      sext1770_2514 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2528_inst
    process(tmp655_2504) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp655_2504, type_cast_2527_wire_constant, tmp_var);
      sext1722_2529 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2552_inst
    process(mul675_2543) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul675_2543, type_cast_2551_wire_constant, tmp_var);
      sext1771_2553 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2567_inst
    process(conv686_2547) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv686_2547, type_cast_2566_wire_constant, tmp_var);
      shl810_2568 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2573_inst
    process(conv664_2508) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv664_2508, type_cast_2572_wire_constant, tmp_var);
      mul667_2574 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3062_inst
    process(tmp867_3041) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp867_3041, type_cast_3061_wire_constant, tmp_var);
      sext1772_3063 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3077_inst
    process(tmp871_3053) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp871_3053, type_cast_3076_wire_constant, tmp_var);
      sext1724_3078 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3101_inst
    process(mul891_3092) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul891_3092, type_cast_3100_wire_constant, tmp_var);
      sext1773_3102 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3116_inst
    process(conv902_3096) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv902_3096, type_cast_3115_wire_constant, tmp_var);
      shl1029_3117 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3122_inst
    process(conv880_3057) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv880_3057, type_cast_3121_wire_constant, tmp_var);
      mul883_3123 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3651_inst
    process(tmp1091_3630) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp1091_3630, type_cast_3650_wire_constant, tmp_var);
      sext1774_3652 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3666_inst
    process(tmp1095_3642) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp1095_3642, type_cast_3665_wire_constant, tmp_var);
      sext1726_3667 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3690_inst
    process(mul1115_3681) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul1115_3681, type_cast_3689_wire_constant, tmp_var);
      sext1775_3691 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3705_inst
    process(conv1126_3685) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1126_3685, type_cast_3704_wire_constant, tmp_var);
      shl1251_3706 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3711_inst
    process(conv1104_3646) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1104_3646, type_cast_3710_wire_constant, tmp_var);
      mul1107_3712 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4218_inst
    process(tmp1310_4197) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp1310_4197, type_cast_4217_wire_constant, tmp_var);
      sext1776_4219 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4233_inst
    process(tmp1314_4209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp1314_4209, type_cast_4232_wire_constant, tmp_var);
      sext1728_4234 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4257_inst
    process(mul1334_4248) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul1334_4248, type_cast_4256_wire_constant, tmp_var);
      sext1777_4258 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4272_inst
    process(conv1345_4252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1345_4252, type_cast_4271_wire_constant, tmp_var);
      shl1470_4273 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4278_inst
    process(conv1323_4213) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1323_4213, type_cast_4277_wire_constant, tmp_var);
      mul1326_4279 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4789_inst
    process(tmp1531_4768) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp1531_4768, type_cast_4788_wire_constant, tmp_var);
      sext1778_4790 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4804_inst
    process(tmp1535_4780) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp1535_4780, type_cast_4803_wire_constant, tmp_var);
      sext1730_4805 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4828_inst
    process(mul1555_4819) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul1555_4819, type_cast_4827_wire_constant, tmp_var);
      sext1779_4829 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4843_inst
    process(conv1566_4823) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1566_4823, type_cast_4842_wire_constant, tmp_var);
      shl1689_4844 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4849_inst
    process(conv1544_4784) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1544_4784, type_cast_4848_wire_constant, tmp_var);
      mul1547_4850 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_820_inst
    process(tmp21_795) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp21_795, type_cast_819_wire_constant, tmp_var);
      sext1764_821 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_836_inst
    process(tmp24_807) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp24_807, type_cast_835_wire_constant, tmp_var);
      sext_837 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_860_inst
    process(mul40_851) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul40_851, type_cast_859_wire_constant, tmp_var);
      sext1765_861 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_875_inst
    process(conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv48_855, type_cast_874_wire_constant, tmp_var);
      shl_876 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_881_inst
    process(conv31_811) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv31_811, type_cast_880_wire_constant, tmp_var);
      mul_882 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1014_inst
    process(type_cast_1011_wire, type_cast_1013_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1011_wire, type_cast_1013_wire, tmp_var);
      cmp74_1015 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1205_inst
    process(type_cast_1202_wire, type_cast_1204_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1202_wire, type_cast_1204_wire, tmp_var);
      cmp143_1206 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1495_inst
    process(type_cast_1492_wire, type_cast_1494_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1492_wire, type_cast_1494_wire, tmp_var);
      cmp249_1496 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1527_inst
    process(type_cast_1524_wire, type_cast_1526_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1524_wire, type_cast_1526_wire, tmp_var);
      cmp260_1528 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1546_inst
    process(type_cast_1543_wire, type_cast_1545_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1543_wire, type_cast_1545_wire, tmp_var);
      cmp267_1547 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1572_inst
    process(type_cast_1569_wire, type_cast_1571_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1569_wire, type_cast_1571_wire, tmp_var);
      cmp277_1573 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1762_inst
    process(type_cast_1759_wire, type_cast_1761_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1759_wire, type_cast_1761_wire, tmp_var);
      cmp356_1763 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2045_inst
    process(type_cast_2042_wire, type_cast_2044_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2042_wire, type_cast_2044_wire, tmp_var);
      cmp465_2046 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2077_inst
    process(type_cast_2074_wire, type_cast_2076_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2074_wire, type_cast_2076_wire, tmp_var);
      cmp476_2078 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2096_inst
    process(type_cast_2093_wire, type_cast_2095_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2093_wire, type_cast_2095_wire, tmp_var);
      cmp483_2097 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2128_inst
    process(type_cast_2125_wire, type_cast_2127_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2125_wire, type_cast_2127_wire, tmp_var);
      cmp494_2129 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2318_inst
    process(type_cast_2315_wire, type_cast_2317_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2315_wire, type_cast_2317_wire, tmp_var);
      cmp573_2319 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2621_inst
    process(type_cast_2618_wire, type_cast_2620_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2618_wire, type_cast_2620_wire, tmp_var);
      cmp687_2622 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2653_inst
    process(type_cast_2650_wire, type_cast_2652_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2650_wire, type_cast_2652_wire, tmp_var);
      cmp698_2654 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2672_inst
    process(type_cast_2669_wire, type_cast_2671_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2669_wire, type_cast_2671_wire, tmp_var);
      cmp705_2673 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2698_inst
    process(type_cast_2695_wire, type_cast_2697_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2695_wire, type_cast_2697_wire, tmp_var);
      cmp715_2699 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2888_inst
    process(type_cast_2885_wire, type_cast_2887_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2885_wire, type_cast_2887_wire, tmp_var);
      cmp794_2889 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3171_inst
    process(type_cast_3168_wire, type_cast_3170_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3168_wire, type_cast_3170_wire, tmp_var);
      cmp903_3172 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3209_inst
    process(type_cast_3206_wire, type_cast_3208_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3206_wire, type_cast_3208_wire, tmp_var);
      cmp915_3210 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3228_inst
    process(type_cast_3225_wire, type_cast_3227_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3225_wire, type_cast_3227_wire, tmp_var);
      cmp922_3229 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3260_inst
    process(type_cast_3257_wire, type_cast_3259_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3257_wire, type_cast_3259_wire, tmp_var);
      cmp933_3261 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3450_inst
    process(type_cast_3447_wire, type_cast_3449_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3447_wire, type_cast_3449_wire, tmp_var);
      cmp1012_3451 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3759_inst
    process(type_cast_3756_wire, type_cast_3758_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3756_wire, type_cast_3758_wire, tmp_var);
      cmp1127_3760 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3797_inst
    process(type_cast_3794_wire, type_cast_3796_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3794_wire, type_cast_3796_wire, tmp_var);
      cmp1139_3798 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3816_inst
    process(type_cast_3813_wire, type_cast_3815_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3813_wire, type_cast_3815_wire, tmp_var);
      cmp1146_3817 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3842_inst
    process(type_cast_3839_wire, type_cast_3841_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3839_wire, type_cast_3841_wire, tmp_var);
      cmp1156_3843 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4032_inst
    process(type_cast_4029_wire, type_cast_4031_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4029_wire, type_cast_4031_wire, tmp_var);
      cmp1235_4033 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4327_inst
    process(type_cast_4324_wire, type_cast_4326_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4324_wire, type_cast_4326_wire, tmp_var);
      cmp1346_4328 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4353_inst
    process(type_cast_4350_wire, type_cast_4352_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4350_wire, type_cast_4352_wire, tmp_var);
      cmp1356_4354 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4372_inst
    process(type_cast_4369_wire, type_cast_4371_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4369_wire, type_cast_4371_wire, tmp_var);
      cmp1363_4373 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4404_inst
    process(type_cast_4401_wire, type_cast_4403_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4401_wire, type_cast_4403_wire, tmp_var);
      cmp1374_4405 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4594_inst
    process(type_cast_4591_wire, type_cast_4593_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4591_wire, type_cast_4593_wire, tmp_var);
      cmp1453_4595 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4897_inst
    process(type_cast_4894_wire, type_cast_4896_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4894_wire, type_cast_4896_wire, tmp_var);
      cmp1567_4898 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4923_inst
    process(type_cast_4920_wire, type_cast_4922_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4920_wire, type_cast_4922_wire, tmp_var);
      cmp1577_4924 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4942_inst
    process(type_cast_4939_wire, type_cast_4941_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4939_wire, type_cast_4941_wire, tmp_var);
      cmp1584_4943 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4968_inst
    process(type_cast_4965_wire, type_cast_4967_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4965_wire, type_cast_4967_wire, tmp_var);
      cmp1594_4969 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_5158_inst
    process(type_cast_5155_wire, type_cast_5157_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_5155_wire, type_cast_5157_wire, tmp_var);
      cmp1673_5159 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_931_inst
    process(type_cast_928_wire, type_cast_930_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_928_wire, type_cast_930_wire, tmp_var);
      cmp_932 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_963_inst
    process(type_cast_960_wire, type_cast_962_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_960_wire, type_cast_962_wire, tmp_var);
      cmp56_964 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_982_inst
    process(type_cast_979_wire, type_cast_981_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_979_wire, type_cast_981_wire, tmp_var);
      cmp63_983 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1090_inst
    process(conv60_976, conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv60_976, conv48_855, tmp_var);
      sub_1091 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1100_inst
    process(conv46_925, conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv46_925, conv48_855, tmp_var);
      sub109_1101 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1647_inst
    process(conv264_1540, conv248_1420) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv264_1540, conv248_1420, tmp_var);
      sub311_1648 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1657_inst
    process(conv246_1489, conv248_1420) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv246_1489, conv248_1420, tmp_var);
      sub320_1658 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2203_inst
    process(conv480_2090, conv464_1970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv480_2090, conv464_1970, tmp_var);
      sub528_2204 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2213_inst
    process(conv462_2039, conv464_1970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv462_2039, conv464_1970, tmp_var);
      sub537_2214 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2773_inst
    process(conv702_2666, conv686_2547) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv702_2666, conv686_2547, tmp_var);
      sub749_2774 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2783_inst
    process(conv684_2615, conv686_2547) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv684_2615, conv686_2547, tmp_var);
      sub758_2784 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3335_inst
    process(conv919_3222, conv902_3096) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv919_3222, conv902_3096, tmp_var);
      sub967_3336 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3345_inst
    process(conv900_3165, conv902_3096) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv900_3165, conv902_3096, tmp_var);
      sub976_3346 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3917_inst
    process(conv1143_3810, conv1126_3685) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1143_3810, conv1126_3685, tmp_var);
      sub1190_3918 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3927_inst
    process(conv1124_3753, conv1126_3685) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1124_3753, conv1126_3685, tmp_var);
      sub1199_3928 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_4479_inst
    process(conv1360_4366, conv1345_4252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1360_4366, conv1345_4252, tmp_var);
      sub1408_4480 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_4489_inst
    process(conv1343_4321, conv1345_4252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1343_4321, conv1345_4252, tmp_var);
      sub1417_4490 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_5043_inst
    process(conv1581_4936, conv1566_4823) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1581_4936, conv1566_4823, tmp_var);
      sub1628_5044 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_5053_inst
    process(conv1564_4891, conv1566_4823) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1564_4891, conv1566_4823, tmp_var);
      sub1637_5054 <= tmp_var; --
    end process;
    -- shared split operator group (380) : array_obj_ref_1072_index_offset 
    ApIntAdd_group_380: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1071_scaled;
      array_obj_ref_1072_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1072_index_offset_req_0;
      array_obj_ref_1072_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1072_index_offset_req_1;
      array_obj_ref_1072_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_380_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_380_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_380",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 380
    -- shared split operator group (381) : array_obj_ref_1155_index_offset 
    ApIntAdd_group_381: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom130_1154_scaled;
      array_obj_ref_1155_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1155_index_offset_req_0;
      array_obj_ref_1155_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1155_index_offset_req_1;
      array_obj_ref_1155_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_381_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_381_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_381",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 381
    -- shared split operator group (382) : array_obj_ref_1180_index_offset 
    ApIntAdd_group_382: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom135_1179_scaled;
      array_obj_ref_1180_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1180_index_offset_req_0;
      array_obj_ref_1180_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1180_index_offset_req_1;
      array_obj_ref_1180_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_382_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_382_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_382",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 382
    -- shared split operator group (383) : array_obj_ref_1629_index_offset 
    ApIntAdd_group_383: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom298_1628_scaled;
      array_obj_ref_1629_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1629_index_offset_req_0;
      array_obj_ref_1629_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1629_index_offset_req_1;
      array_obj_ref_1629_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_383_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_383_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_383",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 383
    -- shared split operator group (384) : array_obj_ref_1712_index_offset 
    ApIntAdd_group_384: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom341_1711_scaled;
      array_obj_ref_1712_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1712_index_offset_req_0;
      array_obj_ref_1712_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1712_index_offset_req_1;
      array_obj_ref_1712_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_384_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_384_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_384",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 384
    -- shared split operator group (385) : array_obj_ref_1737_index_offset 
    ApIntAdd_group_385: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom346_1736_scaled;
      array_obj_ref_1737_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1737_index_offset_req_0;
      array_obj_ref_1737_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1737_index_offset_req_1;
      array_obj_ref_1737_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_385_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_385_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_385",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 385
    -- shared split operator group (386) : array_obj_ref_2185_index_offset 
    ApIntAdd_group_386: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom515_2184_scaled;
      array_obj_ref_2185_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2185_index_offset_req_0;
      array_obj_ref_2185_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2185_index_offset_req_1;
      array_obj_ref_2185_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_386_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_386_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_386",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 386
    -- shared split operator group (387) : array_obj_ref_2268_index_offset 
    ApIntAdd_group_387: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom558_2267_scaled;
      array_obj_ref_2268_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2268_index_offset_req_0;
      array_obj_ref_2268_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2268_index_offset_req_1;
      array_obj_ref_2268_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_387_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_387_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_387",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 387
    -- shared split operator group (388) : array_obj_ref_2293_index_offset 
    ApIntAdd_group_388: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom563_2292_scaled;
      array_obj_ref_2293_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2293_index_offset_req_0;
      array_obj_ref_2293_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2293_index_offset_req_1;
      array_obj_ref_2293_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_388_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_388_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_388",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 388
    -- shared split operator group (389) : array_obj_ref_2755_index_offset 
    ApIntAdd_group_389: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom736_2754_scaled;
      array_obj_ref_2755_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2755_index_offset_req_0;
      array_obj_ref_2755_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2755_index_offset_req_1;
      array_obj_ref_2755_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_389_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_389_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_389",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 389
    -- shared split operator group (390) : array_obj_ref_2838_index_offset 
    ApIntAdd_group_390: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom779_2837_scaled;
      array_obj_ref_2838_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2838_index_offset_req_0;
      array_obj_ref_2838_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2838_index_offset_req_1;
      array_obj_ref_2838_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_390_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_390_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_390",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 390
    -- shared split operator group (391) : array_obj_ref_2863_index_offset 
    ApIntAdd_group_391: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom784_2862_scaled;
      array_obj_ref_2863_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2863_index_offset_req_0;
      array_obj_ref_2863_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2863_index_offset_req_1;
      array_obj_ref_2863_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_391_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_391_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_391",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 391
    -- shared split operator group (392) : array_obj_ref_3317_index_offset 
    ApIntAdd_group_392: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom954_3316_scaled;
      array_obj_ref_3317_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3317_index_offset_req_0;
      array_obj_ref_3317_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3317_index_offset_req_1;
      array_obj_ref_3317_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_392_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_392_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_392",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 392
    -- shared split operator group (393) : array_obj_ref_3400_index_offset 
    ApIntAdd_group_393: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom997_3399_scaled;
      array_obj_ref_3400_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3400_index_offset_req_0;
      array_obj_ref_3400_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3400_index_offset_req_1;
      array_obj_ref_3400_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_393_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_393_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_393",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 393
    -- shared split operator group (394) : array_obj_ref_3425_index_offset 
    ApIntAdd_group_394: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1002_3424_scaled;
      array_obj_ref_3425_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3425_index_offset_req_0;
      array_obj_ref_3425_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3425_index_offset_req_1;
      array_obj_ref_3425_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_394_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_394_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_394",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 394
    -- shared split operator group (395) : array_obj_ref_3899_index_offset 
    ApIntAdd_group_395: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1177_3898_scaled;
      array_obj_ref_3899_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3899_index_offset_req_0;
      array_obj_ref_3899_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3899_index_offset_req_1;
      array_obj_ref_3899_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_395_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_395_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_395",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 395
    -- shared split operator group (396) : array_obj_ref_3982_index_offset 
    ApIntAdd_group_396: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1220_3981_scaled;
      array_obj_ref_3982_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3982_index_offset_req_0;
      array_obj_ref_3982_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3982_index_offset_req_1;
      array_obj_ref_3982_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_396_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_396_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_396",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 396
    -- shared split operator group (397) : array_obj_ref_4007_index_offset 
    ApIntAdd_group_397: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1225_4006_scaled;
      array_obj_ref_4007_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4007_index_offset_req_0;
      array_obj_ref_4007_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4007_index_offset_req_1;
      array_obj_ref_4007_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_397_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_397_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_397",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 397
    -- shared split operator group (398) : array_obj_ref_4461_index_offset 
    ApIntAdd_group_398: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1395_4460_scaled;
      array_obj_ref_4461_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4461_index_offset_req_0;
      array_obj_ref_4461_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4461_index_offset_req_1;
      array_obj_ref_4461_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_398_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_398_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_398",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 398
    -- shared split operator group (399) : array_obj_ref_4544_index_offset 
    ApIntAdd_group_399: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1438_4543_scaled;
      array_obj_ref_4544_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4544_index_offset_req_0;
      array_obj_ref_4544_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4544_index_offset_req_1;
      array_obj_ref_4544_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_399_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_399_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_399",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 399
    -- shared split operator group (400) : array_obj_ref_4569_index_offset 
    ApIntAdd_group_400: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1443_4568_scaled;
      array_obj_ref_4569_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4569_index_offset_req_0;
      array_obj_ref_4569_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4569_index_offset_req_1;
      array_obj_ref_4569_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_400_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_400_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_400",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 400
    -- shared split operator group (401) : array_obj_ref_5025_index_offset 
    ApIntAdd_group_401: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1615_5024_scaled;
      array_obj_ref_5025_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_5025_index_offset_req_0;
      array_obj_ref_5025_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_5025_index_offset_req_1;
      array_obj_ref_5025_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_401_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_401_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_401",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 401
    -- shared split operator group (402) : array_obj_ref_5108_index_offset 
    ApIntAdd_group_402: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1658_5107_scaled;
      array_obj_ref_5108_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_5108_index_offset_req_0;
      array_obj_ref_5108_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_5108_index_offset_req_1;
      array_obj_ref_5108_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_402_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_402_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_402",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 402
    -- shared split operator group (403) : array_obj_ref_5133_index_offset 
    ApIntAdd_group_403: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1663_5132_scaled;
      array_obj_ref_5133_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_5133_index_offset_req_0;
      array_obj_ref_5133_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_5133_index_offset_req_1;
      array_obj_ref_5133_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_403_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_403_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_403",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 403
    -- unary operator type_cast_1025_inst
    process(kx_x1_913) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_913, tmp_var);
      type_cast_1025_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1030_inst
    process(jx_x1_899) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_899, tmp_var);
      type_cast_1030_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1065_inst
    process(shr_1061) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1061, tmp_var);
      type_cast_1065_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1084_inst
    process(kx_x1_913) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_913, tmp_var);
      type_cast_1084_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1148_inst
    process(shr129_1145) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr129_1145, tmp_var);
      type_cast_1148_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1173_inst
    process(shr134_1170) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr134_1170, tmp_var);
      type_cast_1173_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1191_inst
    process(kx_x1_913) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_913, tmp_var);
      type_cast_1191_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1230_inst
    process(inc_1227) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1227, tmp_var);
      type_cast_1230_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1274_inst
    process(inc165x_xix_x2_1264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc165x_xix_x2_1264, tmp_var);
      type_cast_1274_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1487_inst
    process(i194x_x2_1470) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i194x_x2_1470, tmp_var);
      type_cast_1487_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1538_inst
    process(j240x_x1_1464) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j240x_x1_1464, tmp_var);
      type_cast_1538_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1583_inst
    process(k186x_x1_1477) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k186x_x1_1477, tmp_var);
      type_cast_1583_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1588_inst
    process(j240x_x1_1464) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j240x_x1_1464, tmp_var);
      type_cast_1588_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1622_inst
    process(shr297_1619) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr297_1619, tmp_var);
      type_cast_1622_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1641_inst
    process(k186x_x1_1477) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k186x_x1_1477, tmp_var);
      type_cast_1641_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1705_inst
    process(shr340_1702) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr340_1702, tmp_var);
      type_cast_1705_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1730_inst
    process(shr345_1727) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr345_1727, tmp_var);
      type_cast_1730_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1748_inst
    process(k186x_x1_1477) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k186x_x1_1477, tmp_var);
      type_cast_1748_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1787_inst
    process(inc365_1784) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc365_1784, tmp_var);
      type_cast_1787_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1824_inst
    process(inc379x_xi194x_x2_1815) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc379x_xi194x_x2_1815, tmp_var);
      type_cast_1824_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2037_inst
    process(i406x_x2_2021) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i406x_x2_2021, tmp_var);
      type_cast_2037_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2088_inst
    process(j456x_x1_2027) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j456x_x1_2027, tmp_var);
      type_cast_2088_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2139_inst
    process(k402x_x1_2014) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k402x_x1_2014, tmp_var);
      type_cast_2139_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2144_inst
    process(j456x_x1_2027) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j456x_x1_2027, tmp_var);
      type_cast_2144_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2178_inst
    process(shr514_2175) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr514_2175, tmp_var);
      type_cast_2178_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2197_inst
    process(k402x_x1_2014) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k402x_x1_2014, tmp_var);
      type_cast_2197_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2261_inst
    process(shr557_2258) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr557_2258, tmp_var);
      type_cast_2261_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2286_inst
    process(shr562_2283) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr562_2283, tmp_var);
      type_cast_2286_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2304_inst
    process(k402x_x1_2014) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k402x_x1_2014, tmp_var);
      type_cast_2304_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2343_inst
    process(inc582_2340) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc582_2340, tmp_var);
      type_cast_2343_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2387_inst
    process(inc597x_xi406x_x2_2377) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc597x_xi406x_x2_2377, tmp_var);
      type_cast_2387_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2613_inst
    process(i628x_x2_2598) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i628x_x2_2598, tmp_var);
      type_cast_2613_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2664_inst
    process(j678x_x1_2604) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j678x_x1_2604, tmp_var);
      type_cast_2664_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2709_inst
    process(k620x_x1_2591) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k620x_x1_2591, tmp_var);
      type_cast_2709_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2714_inst
    process(j678x_x1_2604) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j678x_x1_2604, tmp_var);
      type_cast_2714_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2748_inst
    process(shr735_2745) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr735_2745, tmp_var);
      type_cast_2748_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2767_inst
    process(k620x_x1_2591) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k620x_x1_2591, tmp_var);
      type_cast_2767_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2831_inst
    process(shr778_2828) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr778_2828, tmp_var);
      type_cast_2831_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2856_inst
    process(shr783_2853) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr783_2853, tmp_var);
      type_cast_2856_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2874_inst
    process(k620x_x1_2591) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k620x_x1_2591, tmp_var);
      type_cast_2874_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2913_inst
    process(inc803_2910) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc803_2910, tmp_var);
      type_cast_2913_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2950_inst
    process(inc817x_xi628x_x2_2941) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc817x_xi628x_x2_2941, tmp_var);
      type_cast_2950_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3163_inst
    process(i844x_x2_3147) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i844x_x2_3147, tmp_var);
      type_cast_3163_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3220_inst
    process(j894x_x1_3153) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j894x_x1_3153, tmp_var);
      type_cast_3220_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3271_inst
    process(k840x_x1_3140) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k840x_x1_3140, tmp_var);
      type_cast_3271_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3276_inst
    process(j894x_x1_3153) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j894x_x1_3153, tmp_var);
      type_cast_3276_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3310_inst
    process(shr953_3307) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr953_3307, tmp_var);
      type_cast_3310_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3329_inst
    process(k840x_x1_3140) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k840x_x1_3140, tmp_var);
      type_cast_3329_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3393_inst
    process(shr996_3390) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr996_3390, tmp_var);
      type_cast_3393_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3418_inst
    process(shr1001_3415) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1001_3415, tmp_var);
      type_cast_3418_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3436_inst
    process(k840x_x1_3140) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k840x_x1_3140, tmp_var);
      type_cast_3436_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3475_inst
    process(inc1021_3472) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1021_3472, tmp_var);
      type_cast_3475_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3519_inst
    process(inc1036x_xi844x_x2_3509) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1036x_xi844x_x2_3509, tmp_var);
      type_cast_3519_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3751_inst
    process(i1068x_x2_3736) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i1068x_x2_3736, tmp_var);
      type_cast_3751_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3808_inst
    process(j1118x_x1_3742) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1118x_x1_3742, tmp_var);
      type_cast_3808_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3853_inst
    process(k1060x_x1_3729) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1060x_x1_3729, tmp_var);
      type_cast_3853_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3858_inst
    process(j1118x_x1_3742) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1118x_x1_3742, tmp_var);
      type_cast_3858_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3892_inst
    process(shr1176_3889) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1176_3889, tmp_var);
      type_cast_3892_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3911_inst
    process(k1060x_x1_3729) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1060x_x1_3729, tmp_var);
      type_cast_3911_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3975_inst
    process(shr1219_3972) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1219_3972, tmp_var);
      type_cast_3975_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4000_inst
    process(shr1224_3997) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1224_3997, tmp_var);
      type_cast_4000_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4018_inst
    process(k1060x_x1_3729) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1060x_x1_3729, tmp_var);
      type_cast_4018_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4057_inst
    process(inc1244_4054) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1244_4054, tmp_var);
      type_cast_4057_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4094_inst
    process(inc1258x_xi1068x_x2_4085) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1258x_xi1068x_x2_4085, tmp_var);
      type_cast_4094_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4319_inst
    process(i1286x_x2_4303) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i1286x_x2_4303, tmp_var);
      type_cast_4319_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4364_inst
    process(j1337x_x1_4309) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1337x_x1_4309, tmp_var);
      type_cast_4364_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4415_inst
    process(k1282x_x1_4296) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1282x_x1_4296, tmp_var);
      type_cast_4415_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4420_inst
    process(j1337x_x1_4309) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1337x_x1_4309, tmp_var);
      type_cast_4420_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4454_inst
    process(shr1394_4451) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1394_4451, tmp_var);
      type_cast_4454_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4473_inst
    process(k1282x_x1_4296) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1282x_x1_4296, tmp_var);
      type_cast_4473_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4537_inst
    process(shr1437_4534) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1437_4534, tmp_var);
      type_cast_4537_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4562_inst
    process(shr1442_4559) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1442_4559, tmp_var);
      type_cast_4562_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4580_inst
    process(k1282x_x1_4296) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1282x_x1_4296, tmp_var);
      type_cast_4580_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4619_inst
    process(inc1462_4616) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1462_4616, tmp_var);
      type_cast_4619_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4663_inst
    process(inc1477x_xi1286x_x2_4653) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1477x_xi1286x_x2_4653, tmp_var);
      type_cast_4663_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4889_inst
    process(i1507x_x2_4874) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i1507x_x2_4874, tmp_var);
      type_cast_4889_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4934_inst
    process(j1558x_x1_4880) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1558x_x1_4880, tmp_var);
      type_cast_4934_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4979_inst
    process(k1499x_x1_4867) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1499x_x1_4867, tmp_var);
      type_cast_4979_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4984_inst
    process(j1558x_x1_4880) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1558x_x1_4880, tmp_var);
      type_cast_4984_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5018_inst
    process(shr1614_5015) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1614_5015, tmp_var);
      type_cast_5018_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5037_inst
    process(k1499x_x1_4867) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1499x_x1_4867, tmp_var);
      type_cast_5037_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5101_inst
    process(shr1657_5098) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1657_5098, tmp_var);
      type_cast_5101_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5126_inst
    process(shr1662_5123) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1662_5123, tmp_var);
      type_cast_5126_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5144_inst
    process(k1499x_x1_4867) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1499x_x1_4867, tmp_var);
      type_cast_5144_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5183_inst
    process(inc1682_5180) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1682_5180, tmp_var);
      type_cast_5183_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5220_inst
    process(inc1696x_xi1507x_x2_5211) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1696x_xi1507x_x2_5211, tmp_var);
      type_cast_5220_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_923_inst
    process(ix_x2_906) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_906, tmp_var);
      type_cast_923_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_974_inst
    process(jx_x1_899) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_899, tmp_var);
      type_cast_974_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_col_high_992_load_0 LOAD_col_high_782_load_0 LOAD_col_high_1791_load_0 LOAD_col_high_1234_load_0 LOAD_col_high_4061_load_0 LOAD_col_high_3238_load_0 LOAD_col_high_2106_load_0 LOAD_col_high_1556_load_0 LOAD_col_high_2347_load_0 LOAD_col_high_4382_load_0 LOAD_col_high_2682_load_0 LOAD_col_high_2917_load_0 LOAD_col_high_3479_load_0 LOAD_col_high_5187_load_0 LOAD_col_high_3826_load_0 LOAD_col_high_4623_load_0 LOAD_col_high_4952_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(16 downto 0);
      signal data_out: std_logic_vector(135 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 16 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 16 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 16 downto 0);
      signal guard_vector : std_logic_vector( 16 downto 0);
      constant inBUFs : IntegerArray(16 downto 0) := (16 => 0, 15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(16 downto 0) := (16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(16 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false);
      constant guardBuffering: IntegerArray(16 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2);
      -- 
    begin -- 
      reqL_unguarded(16) <= LOAD_col_high_992_load_0_req_0;
      reqL_unguarded(15) <= LOAD_col_high_782_load_0_req_0;
      reqL_unguarded(14) <= LOAD_col_high_1791_load_0_req_0;
      reqL_unguarded(13) <= LOAD_col_high_1234_load_0_req_0;
      reqL_unguarded(12) <= LOAD_col_high_4061_load_0_req_0;
      reqL_unguarded(11) <= LOAD_col_high_3238_load_0_req_0;
      reqL_unguarded(10) <= LOAD_col_high_2106_load_0_req_0;
      reqL_unguarded(9) <= LOAD_col_high_1556_load_0_req_0;
      reqL_unguarded(8) <= LOAD_col_high_2347_load_0_req_0;
      reqL_unguarded(7) <= LOAD_col_high_4382_load_0_req_0;
      reqL_unguarded(6) <= LOAD_col_high_2682_load_0_req_0;
      reqL_unguarded(5) <= LOAD_col_high_2917_load_0_req_0;
      reqL_unguarded(4) <= LOAD_col_high_3479_load_0_req_0;
      reqL_unguarded(3) <= LOAD_col_high_5187_load_0_req_0;
      reqL_unguarded(2) <= LOAD_col_high_3826_load_0_req_0;
      reqL_unguarded(1) <= LOAD_col_high_4623_load_0_req_0;
      reqL_unguarded(0) <= LOAD_col_high_4952_load_0_req_0;
      LOAD_col_high_992_load_0_ack_0 <= ackL_unguarded(16);
      LOAD_col_high_782_load_0_ack_0 <= ackL_unguarded(15);
      LOAD_col_high_1791_load_0_ack_0 <= ackL_unguarded(14);
      LOAD_col_high_1234_load_0_ack_0 <= ackL_unguarded(13);
      LOAD_col_high_4061_load_0_ack_0 <= ackL_unguarded(12);
      LOAD_col_high_3238_load_0_ack_0 <= ackL_unguarded(11);
      LOAD_col_high_2106_load_0_ack_0 <= ackL_unguarded(10);
      LOAD_col_high_1556_load_0_ack_0 <= ackL_unguarded(9);
      LOAD_col_high_2347_load_0_ack_0 <= ackL_unguarded(8);
      LOAD_col_high_4382_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_col_high_2682_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_col_high_2917_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_col_high_3479_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_col_high_5187_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_col_high_3826_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_col_high_4623_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_col_high_4952_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(16) <= LOAD_col_high_992_load_0_req_1;
      reqR_unguarded(15) <= LOAD_col_high_782_load_0_req_1;
      reqR_unguarded(14) <= LOAD_col_high_1791_load_0_req_1;
      reqR_unguarded(13) <= LOAD_col_high_1234_load_0_req_1;
      reqR_unguarded(12) <= LOAD_col_high_4061_load_0_req_1;
      reqR_unguarded(11) <= LOAD_col_high_3238_load_0_req_1;
      reqR_unguarded(10) <= LOAD_col_high_2106_load_0_req_1;
      reqR_unguarded(9) <= LOAD_col_high_1556_load_0_req_1;
      reqR_unguarded(8) <= LOAD_col_high_2347_load_0_req_1;
      reqR_unguarded(7) <= LOAD_col_high_4382_load_0_req_1;
      reqR_unguarded(6) <= LOAD_col_high_2682_load_0_req_1;
      reqR_unguarded(5) <= LOAD_col_high_2917_load_0_req_1;
      reqR_unguarded(4) <= LOAD_col_high_3479_load_0_req_1;
      reqR_unguarded(3) <= LOAD_col_high_5187_load_0_req_1;
      reqR_unguarded(2) <= LOAD_col_high_3826_load_0_req_1;
      reqR_unguarded(1) <= LOAD_col_high_4623_load_0_req_1;
      reqR_unguarded(0) <= LOAD_col_high_4952_load_0_req_1;
      LOAD_col_high_992_load_0_ack_1 <= ackR_unguarded(16);
      LOAD_col_high_782_load_0_ack_1 <= ackR_unguarded(15);
      LOAD_col_high_1791_load_0_ack_1 <= ackR_unguarded(14);
      LOAD_col_high_1234_load_0_ack_1 <= ackR_unguarded(13);
      LOAD_col_high_4061_load_0_ack_1 <= ackR_unguarded(12);
      LOAD_col_high_3238_load_0_ack_1 <= ackR_unguarded(11);
      LOAD_col_high_2106_load_0_ack_1 <= ackR_unguarded(10);
      LOAD_col_high_1556_load_0_ack_1 <= ackR_unguarded(9);
      LOAD_col_high_2347_load_0_ack_1 <= ackR_unguarded(8);
      LOAD_col_high_4382_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_col_high_2682_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_col_high_2917_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_col_high_3479_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_col_high_5187_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_col_high_3826_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_col_high_4623_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_col_high_4952_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_15: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_16: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_16", num_slots => 1) -- 
        port map (req => reqL_unregulated(16), -- 
          ack => ackL_unregulated(16),
          regulated_req => reqL(16),
          regulated_ack => ackL(16),
          release_req => reqR(16),
          release_ack => ackR(16),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 17, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_col_high_992_word_address_0 & LOAD_col_high_782_word_address_0 & LOAD_col_high_1791_word_address_0 & LOAD_col_high_1234_word_address_0 & LOAD_col_high_4061_word_address_0 & LOAD_col_high_3238_word_address_0 & LOAD_col_high_2106_word_address_0 & LOAD_col_high_1556_word_address_0 & LOAD_col_high_2347_word_address_0 & LOAD_col_high_4382_word_address_0 & LOAD_col_high_2682_word_address_0 & LOAD_col_high_2917_word_address_0 & LOAD_col_high_3479_word_address_0 & LOAD_col_high_5187_word_address_0 & LOAD_col_high_3826_word_address_0 & LOAD_col_high_4623_word_address_0 & LOAD_col_high_4952_word_address_0;
      LOAD_col_high_992_data_0 <= data_out(135 downto 128);
      LOAD_col_high_782_data_0 <= data_out(127 downto 120);
      LOAD_col_high_1791_data_0 <= data_out(119 downto 112);
      LOAD_col_high_1234_data_0 <= data_out(111 downto 104);
      LOAD_col_high_4061_data_0 <= data_out(103 downto 96);
      LOAD_col_high_3238_data_0 <= data_out(95 downto 88);
      LOAD_col_high_2106_data_0 <= data_out(87 downto 80);
      LOAD_col_high_1556_data_0 <= data_out(79 downto 72);
      LOAD_col_high_2347_data_0 <= data_out(71 downto 64);
      LOAD_col_high_4382_data_0 <= data_out(63 downto 56);
      LOAD_col_high_2682_data_0 <= data_out(55 downto 48);
      LOAD_col_high_2917_data_0 <= data_out(47 downto 40);
      LOAD_col_high_3479_data_0 <= data_out(39 downto 32);
      LOAD_col_high_5187_data_0 <= data_out(31 downto 24);
      LOAD_col_high_3826_data_0 <= data_out(23 downto 16);
      LOAD_col_high_4623_data_0 <= data_out(15 downto 8);
      LOAD_col_high_4952_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 17,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 17,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(7 downto 0),
          mtag => memory_space_2_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : LOAD_depth_high_779_load_0 LOAD_depth_high_1902_load_0 LOAD_depth_high_1352_load_0 LOAD_depth_high_4184_load_0 LOAD_depth_high_2479_load_0 LOAD_depth_high_3028_load_0 LOAD_depth_high_3617_load_0 LOAD_depth_high_4755_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= LOAD_depth_high_779_load_0_req_0;
      reqL_unguarded(6) <= LOAD_depth_high_1902_load_0_req_0;
      reqL_unguarded(5) <= LOAD_depth_high_1352_load_0_req_0;
      reqL_unguarded(4) <= LOAD_depth_high_4184_load_0_req_0;
      reqL_unguarded(3) <= LOAD_depth_high_2479_load_0_req_0;
      reqL_unguarded(2) <= LOAD_depth_high_3028_load_0_req_0;
      reqL_unguarded(1) <= LOAD_depth_high_3617_load_0_req_0;
      reqL_unguarded(0) <= LOAD_depth_high_4755_load_0_req_0;
      LOAD_depth_high_779_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_depth_high_1902_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_depth_high_1352_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_depth_high_4184_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_depth_high_2479_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_depth_high_3028_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_depth_high_3617_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_depth_high_4755_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= LOAD_depth_high_779_load_0_req_1;
      reqR_unguarded(6) <= LOAD_depth_high_1902_load_0_req_1;
      reqR_unguarded(5) <= LOAD_depth_high_1352_load_0_req_1;
      reqR_unguarded(4) <= LOAD_depth_high_4184_load_0_req_1;
      reqR_unguarded(3) <= LOAD_depth_high_2479_load_0_req_1;
      reqR_unguarded(2) <= LOAD_depth_high_3028_load_0_req_1;
      reqR_unguarded(1) <= LOAD_depth_high_3617_load_0_req_1;
      reqR_unguarded(0) <= LOAD_depth_high_4755_load_0_req_1;
      LOAD_depth_high_779_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_depth_high_1902_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_depth_high_1352_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_depth_high_4184_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_depth_high_2479_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_depth_high_3028_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_depth_high_3617_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_depth_high_4755_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_depth_high_779_word_address_0 & LOAD_depth_high_1902_word_address_0 & LOAD_depth_high_1352_word_address_0 & LOAD_depth_high_4184_word_address_0 & LOAD_depth_high_2479_word_address_0 & LOAD_depth_high_3028_word_address_0 & LOAD_depth_high_3617_word_address_0 & LOAD_depth_high_4755_word_address_0;
      LOAD_depth_high_779_data_0 <= data_out(63 downto 56);
      LOAD_depth_high_1902_data_0 <= data_out(55 downto 48);
      LOAD_depth_high_1352_data_0 <= data_out(47 downto 40);
      LOAD_depth_high_4184_data_0 <= data_out(39 downto 32);
      LOAD_depth_high_2479_data_0 <= data_out(31 downto 24);
      LOAD_depth_high_3028_data_0 <= data_out(23 downto 16);
      LOAD_depth_high_3617_data_0 <= data_out(15 downto 8);
      LOAD_depth_high_4755_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 1,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(0 downto 0),
          mtag => memory_space_4_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(7 downto 0),
          mtag => memory_space_4_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : LOAD_pad_776_load_0 LOAD_pad_4181_load_0 LOAD_pad_1899_load_0 LOAD_pad_1349_load_0 LOAD_pad_2476_load_0 LOAD_pad_3025_load_0 LOAD_pad_3614_load_0 LOAD_pad_4752_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= LOAD_pad_776_load_0_req_0;
      reqL_unguarded(6) <= LOAD_pad_4181_load_0_req_0;
      reqL_unguarded(5) <= LOAD_pad_1899_load_0_req_0;
      reqL_unguarded(4) <= LOAD_pad_1349_load_0_req_0;
      reqL_unguarded(3) <= LOAD_pad_2476_load_0_req_0;
      reqL_unguarded(2) <= LOAD_pad_3025_load_0_req_0;
      reqL_unguarded(1) <= LOAD_pad_3614_load_0_req_0;
      reqL_unguarded(0) <= LOAD_pad_4752_load_0_req_0;
      LOAD_pad_776_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_pad_4181_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_pad_1899_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_pad_1349_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_pad_2476_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_pad_3025_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_pad_3614_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_pad_4752_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= LOAD_pad_776_load_0_req_1;
      reqR_unguarded(6) <= LOAD_pad_4181_load_0_req_1;
      reqR_unguarded(5) <= LOAD_pad_1899_load_0_req_1;
      reqR_unguarded(4) <= LOAD_pad_1349_load_0_req_1;
      reqR_unguarded(3) <= LOAD_pad_2476_load_0_req_1;
      reqR_unguarded(2) <= LOAD_pad_3025_load_0_req_1;
      reqR_unguarded(1) <= LOAD_pad_3614_load_0_req_1;
      reqR_unguarded(0) <= LOAD_pad_4752_load_0_req_1;
      LOAD_pad_776_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_pad_4181_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_pad_1899_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_pad_1349_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_pad_2476_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_pad_3025_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_pad_3614_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_pad_4752_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_pad_776_word_address_0 & LOAD_pad_4181_word_address_0 & LOAD_pad_1899_word_address_0 & LOAD_pad_1349_word_address_0 & LOAD_pad_2476_word_address_0 & LOAD_pad_3025_word_address_0 & LOAD_pad_3614_word_address_0 & LOAD_pad_4752_word_address_0;
      LOAD_pad_776_data_0 <= data_out(63 downto 56);
      LOAD_pad_4181_data_0 <= data_out(55 downto 48);
      LOAD_pad_1899_data_0 <= data_out(47 downto 40);
      LOAD_pad_1349_data_0 <= data_out(39 downto 32);
      LOAD_pad_2476_data_0 <= data_out(31 downto 24);
      LOAD_pad_3025_data_0 <= data_out(23 downto 16);
      LOAD_pad_3614_data_0 <= data_out(15 downto 8);
      LOAD_pad_4752_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(7 downto 0),
          mtag => memory_space_7_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : LOAD_row_high_3181_load_0 LOAD_row_high_941_load_0 LOAD_row_high_1828_load_0 LOAD_row_high_1278_load_0 LOAD_row_high_1505_load_0 LOAD_row_high_2055_load_0 LOAD_row_high_4098_load_0 LOAD_row_high_2391_load_0 LOAD_row_high_4337_load_0 LOAD_row_high_2631_load_0 LOAD_row_high_2954_load_0 LOAD_row_high_3523_load_0 LOAD_row_high_3769_load_0 LOAD_row_high_5224_load_0 LOAD_row_high_4667_load_0 LOAD_row_high_4907_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      reqL_unguarded(15) <= LOAD_row_high_3181_load_0_req_0;
      reqL_unguarded(14) <= LOAD_row_high_941_load_0_req_0;
      reqL_unguarded(13) <= LOAD_row_high_1828_load_0_req_0;
      reqL_unguarded(12) <= LOAD_row_high_1278_load_0_req_0;
      reqL_unguarded(11) <= LOAD_row_high_1505_load_0_req_0;
      reqL_unguarded(10) <= LOAD_row_high_2055_load_0_req_0;
      reqL_unguarded(9) <= LOAD_row_high_4098_load_0_req_0;
      reqL_unguarded(8) <= LOAD_row_high_2391_load_0_req_0;
      reqL_unguarded(7) <= LOAD_row_high_4337_load_0_req_0;
      reqL_unguarded(6) <= LOAD_row_high_2631_load_0_req_0;
      reqL_unguarded(5) <= LOAD_row_high_2954_load_0_req_0;
      reqL_unguarded(4) <= LOAD_row_high_3523_load_0_req_0;
      reqL_unguarded(3) <= LOAD_row_high_3769_load_0_req_0;
      reqL_unguarded(2) <= LOAD_row_high_5224_load_0_req_0;
      reqL_unguarded(1) <= LOAD_row_high_4667_load_0_req_0;
      reqL_unguarded(0) <= LOAD_row_high_4907_load_0_req_0;
      LOAD_row_high_3181_load_0_ack_0 <= ackL_unguarded(15);
      LOAD_row_high_941_load_0_ack_0 <= ackL_unguarded(14);
      LOAD_row_high_1828_load_0_ack_0 <= ackL_unguarded(13);
      LOAD_row_high_1278_load_0_ack_0 <= ackL_unguarded(12);
      LOAD_row_high_1505_load_0_ack_0 <= ackL_unguarded(11);
      LOAD_row_high_2055_load_0_ack_0 <= ackL_unguarded(10);
      LOAD_row_high_4098_load_0_ack_0 <= ackL_unguarded(9);
      LOAD_row_high_2391_load_0_ack_0 <= ackL_unguarded(8);
      LOAD_row_high_4337_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_row_high_2631_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_row_high_2954_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_row_high_3523_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_row_high_3769_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_row_high_5224_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_row_high_4667_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_row_high_4907_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= LOAD_row_high_3181_load_0_req_1;
      reqR_unguarded(14) <= LOAD_row_high_941_load_0_req_1;
      reqR_unguarded(13) <= LOAD_row_high_1828_load_0_req_1;
      reqR_unguarded(12) <= LOAD_row_high_1278_load_0_req_1;
      reqR_unguarded(11) <= LOAD_row_high_1505_load_0_req_1;
      reqR_unguarded(10) <= LOAD_row_high_2055_load_0_req_1;
      reqR_unguarded(9) <= LOAD_row_high_4098_load_0_req_1;
      reqR_unguarded(8) <= LOAD_row_high_2391_load_0_req_1;
      reqR_unguarded(7) <= LOAD_row_high_4337_load_0_req_1;
      reqR_unguarded(6) <= LOAD_row_high_2631_load_0_req_1;
      reqR_unguarded(5) <= LOAD_row_high_2954_load_0_req_1;
      reqR_unguarded(4) <= LOAD_row_high_3523_load_0_req_1;
      reqR_unguarded(3) <= LOAD_row_high_3769_load_0_req_1;
      reqR_unguarded(2) <= LOAD_row_high_5224_load_0_req_1;
      reqR_unguarded(1) <= LOAD_row_high_4667_load_0_req_1;
      reqR_unguarded(0) <= LOAD_row_high_4907_load_0_req_1;
      LOAD_row_high_3181_load_0_ack_1 <= ackR_unguarded(15);
      LOAD_row_high_941_load_0_ack_1 <= ackR_unguarded(14);
      LOAD_row_high_1828_load_0_ack_1 <= ackR_unguarded(13);
      LOAD_row_high_1278_load_0_ack_1 <= ackR_unguarded(12);
      LOAD_row_high_1505_load_0_ack_1 <= ackR_unguarded(11);
      LOAD_row_high_2055_load_0_ack_1 <= ackR_unguarded(10);
      LOAD_row_high_4098_load_0_ack_1 <= ackR_unguarded(9);
      LOAD_row_high_2391_load_0_ack_1 <= ackR_unguarded(8);
      LOAD_row_high_4337_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_row_high_2631_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_row_high_2954_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_row_high_3523_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_row_high_3769_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_row_high_5224_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_row_high_4667_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_row_high_4907_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_15: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_row_high_3181_word_address_0 & LOAD_row_high_941_word_address_0 & LOAD_row_high_1828_word_address_0 & LOAD_row_high_1278_word_address_0 & LOAD_row_high_1505_word_address_0 & LOAD_row_high_2055_word_address_0 & LOAD_row_high_4098_word_address_0 & LOAD_row_high_2391_word_address_0 & LOAD_row_high_4337_word_address_0 & LOAD_row_high_2631_word_address_0 & LOAD_row_high_2954_word_address_0 & LOAD_row_high_3523_word_address_0 & LOAD_row_high_3769_word_address_0 & LOAD_row_high_5224_word_address_0 & LOAD_row_high_4667_word_address_0 & LOAD_row_high_4907_word_address_0;
      LOAD_row_high_3181_data_0 <= data_out(127 downto 120);
      LOAD_row_high_941_data_0 <= data_out(119 downto 112);
      LOAD_row_high_1828_data_0 <= data_out(111 downto 104);
      LOAD_row_high_1278_data_0 <= data_out(103 downto 96);
      LOAD_row_high_1505_data_0 <= data_out(95 downto 88);
      LOAD_row_high_2055_data_0 <= data_out(87 downto 80);
      LOAD_row_high_4098_data_0 <= data_out(79 downto 72);
      LOAD_row_high_2391_data_0 <= data_out(71 downto 64);
      LOAD_row_high_4337_data_0 <= data_out(63 downto 56);
      LOAD_row_high_2631_data_0 <= data_out(55 downto 48);
      LOAD_row_high_2954_data_0 <= data_out(47 downto 40);
      LOAD_row_high_3523_data_0 <= data_out(39 downto 32);
      LOAD_row_high_3769_data_0 <= data_out(31 downto 24);
      LOAD_row_high_5224_data_0 <= data_out(23 downto 16);
      LOAD_row_high_4667_data_0 <= data_out(15 downto 8);
      LOAD_row_high_4907_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 1,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 8,
        num_reqs => 16,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(7 downto 0),
          mtag => memory_space_8_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1717_load_0 ptr_deref_1160_load_0 ptr_deref_2273_load_0 ptr_deref_3987_load_0 ptr_deref_2843_load_0 ptr_deref_3405_load_0 ptr_deref_4549_load_0 ptr_deref_5113_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(111 downto 0);
      signal data_out: std_logic_vector(511 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= ptr_deref_1717_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_1160_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_2273_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_3987_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_2843_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_3405_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_4549_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_5113_load_0_req_0;
      ptr_deref_1717_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_1160_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_2273_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_3987_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_2843_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_3405_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_4549_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_5113_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ptr_deref_1717_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_1160_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_2273_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_3987_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_2843_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_3405_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_4549_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_5113_load_0_req_1;
      ptr_deref_1717_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_1160_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_2273_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_3987_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_2843_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_3405_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_4549_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_5113_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1717_word_address_0 & ptr_deref_1160_word_address_0 & ptr_deref_2273_word_address_0 & ptr_deref_3987_word_address_0 & ptr_deref_2843_word_address_0 & ptr_deref_3405_word_address_0 & ptr_deref_4549_word_address_0 & ptr_deref_5113_word_address_0;
      ptr_deref_1717_data_0 <= data_out(511 downto 448);
      ptr_deref_1160_data_0 <= data_out(447 downto 384);
      ptr_deref_2273_data_0 <= data_out(383 downto 320);
      ptr_deref_3987_data_0 <= data_out(319 downto 256);
      ptr_deref_2843_data_0 <= data_out(255 downto 192);
      ptr_deref_3405_data_0 <= data_out(191 downto 128);
      ptr_deref_4549_data_0 <= data_out(127 downto 64);
      ptr_deref_5113_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 14,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 64,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_806_load_0 ptr_deref_794_load_0 ptr_deref_1926_load_0 ptr_deref_1914_load_0 ptr_deref_3052_load_0 ptr_deref_1364_load_0 ptr_deref_1376_load_0 ptr_deref_4196_load_0 ptr_deref_3040_load_0 ptr_deref_4208_load_0 ptr_deref_2491_load_0 ptr_deref_2503_load_0 ptr_deref_3629_load_0 ptr_deref_3641_load_0 ptr_deref_4767_load_0 ptr_deref_4779_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(111 downto 0);
      signal data_out: std_logic_vector(511 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      reqL_unguarded(15) <= ptr_deref_806_load_0_req_0;
      reqL_unguarded(14) <= ptr_deref_794_load_0_req_0;
      reqL_unguarded(13) <= ptr_deref_1926_load_0_req_0;
      reqL_unguarded(12) <= ptr_deref_1914_load_0_req_0;
      reqL_unguarded(11) <= ptr_deref_3052_load_0_req_0;
      reqL_unguarded(10) <= ptr_deref_1364_load_0_req_0;
      reqL_unguarded(9) <= ptr_deref_1376_load_0_req_0;
      reqL_unguarded(8) <= ptr_deref_4196_load_0_req_0;
      reqL_unguarded(7) <= ptr_deref_3040_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_4208_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_2491_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_2503_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_3629_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_3641_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_4767_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_4779_load_0_req_0;
      ptr_deref_806_load_0_ack_0 <= ackL_unguarded(15);
      ptr_deref_794_load_0_ack_0 <= ackL_unguarded(14);
      ptr_deref_1926_load_0_ack_0 <= ackL_unguarded(13);
      ptr_deref_1914_load_0_ack_0 <= ackL_unguarded(12);
      ptr_deref_3052_load_0_ack_0 <= ackL_unguarded(11);
      ptr_deref_1364_load_0_ack_0 <= ackL_unguarded(10);
      ptr_deref_1376_load_0_ack_0 <= ackL_unguarded(9);
      ptr_deref_4196_load_0_ack_0 <= ackL_unguarded(8);
      ptr_deref_3040_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_4208_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_2491_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_2503_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_3629_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_3641_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_4767_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_4779_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= ptr_deref_806_load_0_req_1;
      reqR_unguarded(14) <= ptr_deref_794_load_0_req_1;
      reqR_unguarded(13) <= ptr_deref_1926_load_0_req_1;
      reqR_unguarded(12) <= ptr_deref_1914_load_0_req_1;
      reqR_unguarded(11) <= ptr_deref_3052_load_0_req_1;
      reqR_unguarded(10) <= ptr_deref_1364_load_0_req_1;
      reqR_unguarded(9) <= ptr_deref_1376_load_0_req_1;
      reqR_unguarded(8) <= ptr_deref_4196_load_0_req_1;
      reqR_unguarded(7) <= ptr_deref_3040_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_4208_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_2491_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_2503_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_3629_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_3641_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_4767_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_4779_load_0_req_1;
      ptr_deref_806_load_0_ack_1 <= ackR_unguarded(15);
      ptr_deref_794_load_0_ack_1 <= ackR_unguarded(14);
      ptr_deref_1926_load_0_ack_1 <= ackR_unguarded(13);
      ptr_deref_1914_load_0_ack_1 <= ackR_unguarded(12);
      ptr_deref_3052_load_0_ack_1 <= ackR_unguarded(11);
      ptr_deref_1364_load_0_ack_1 <= ackR_unguarded(10);
      ptr_deref_1376_load_0_ack_1 <= ackR_unguarded(9);
      ptr_deref_4196_load_0_ack_1 <= ackR_unguarded(8);
      ptr_deref_3040_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_4208_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_2491_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_2503_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_3629_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_3641_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_4767_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_4779_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      LoadGroup5_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_15: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_806_word_address_0 & ptr_deref_794_word_address_0 & ptr_deref_1926_word_address_0 & ptr_deref_1914_word_address_0 & ptr_deref_3052_word_address_0 & ptr_deref_1364_word_address_0 & ptr_deref_1376_word_address_0 & ptr_deref_4196_word_address_0 & ptr_deref_3040_word_address_0 & ptr_deref_4208_word_address_0 & ptr_deref_2491_word_address_0 & ptr_deref_2503_word_address_0 & ptr_deref_3629_word_address_0 & ptr_deref_3641_word_address_0 & ptr_deref_4767_word_address_0 & ptr_deref_4779_word_address_0;
      ptr_deref_806_data_0 <= data_out(511 downto 480);
      ptr_deref_794_data_0 <= data_out(479 downto 448);
      ptr_deref_1926_data_0 <= data_out(447 downto 416);
      ptr_deref_1914_data_0 <= data_out(415 downto 384);
      ptr_deref_3052_data_0 <= data_out(383 downto 352);
      ptr_deref_1364_data_0 <= data_out(351 downto 320);
      ptr_deref_1376_data_0 <= data_out(319 downto 288);
      ptr_deref_4196_data_0 <= data_out(287 downto 256);
      ptr_deref_3040_data_0 <= data_out(255 downto 224);
      ptr_deref_4208_data_0 <= data_out(223 downto 192);
      ptr_deref_2491_data_0 <= data_out(191 downto 160);
      ptr_deref_2503_data_0 <= data_out(159 downto 128);
      ptr_deref_3629_data_0 <= data_out(127 downto 96);
      ptr_deref_3641_data_0 <= data_out(95 downto 64);
      ptr_deref_4767_data_0 <= data_out(63 downto 32);
      ptr_deref_4779_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 7,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(6 downto 0),
          mtag => memory_space_6_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 32,
        num_reqs => 16,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(31 downto 0),
          mtag => memory_space_6_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : ptr_deref_746_load_0 ptr_deref_765_load_0 ptr_deref_727_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_746_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_765_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_727_load_0_req_0;
      ptr_deref_746_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_765_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_727_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_746_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_765_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_727_load_0_req_1;
      ptr_deref_746_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_765_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_727_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup6_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup6_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup6_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup6_gI: SplitGuardInterface generic map(name => "LoadGroup6_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_746_word_address_0 & ptr_deref_765_word_address_0 & ptr_deref_727_word_address_0;
      ptr_deref_746_data_0 <= data_out(95 downto 64);
      ptr_deref_765_data_0 <= data_out(63 downto 32);
      ptr_deref_727_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup6", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(6 downto 0),
          mtag => memory_space_5_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup6 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(31 downto 0),
          mtag => memory_space_5_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared store operator group (0) : STORE_col_high_752_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_col_high_752_store_0_req_0;
      STORE_col_high_752_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_col_high_752_store_0_req_1;
      STORE_col_high_752_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_col_high_752_word_address_0;
      data_in <= STORE_col_high_752_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(7 downto 0),
          mtag => memory_space_2_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : STORE_depth_high_771_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_depth_high_771_store_0_req_0;
      STORE_depth_high_771_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_depth_high_771_store_0_req_1;
      STORE_depth_high_771_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_depth_high_771_word_address_0;
      data_in <= STORE_depth_high_771_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(0 downto 0),
          mdata => memory_space_4_sr_data(7 downto 0),
          mtag => memory_space_4_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : STORE_row_high_733_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_row_high_733_store_0_req_0;
      STORE_row_high_733_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_row_high_733_store_0_req_1;
      STORE_row_high_733_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_row_high_733_word_address_0;
      data_in <= STORE_row_high_733_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(7 downto 0),
          mtag => memory_space_8_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_1741_store_0 ptr_deref_1076_store_0 ptr_deref_1184_store_0 ptr_deref_3321_store_0 ptr_deref_1633_store_0 ptr_deref_2189_store_0 ptr_deref_4465_store_0 ptr_deref_2297_store_0 ptr_deref_4011_store_0 ptr_deref_2759_store_0 ptr_deref_2867_store_0 ptr_deref_3429_store_0 ptr_deref_5029_store_0 ptr_deref_5137_store_0 ptr_deref_3903_store_0 ptr_deref_4573_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(223 downto 0);
      signal data_in: std_logic_vector(1023 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      reqL_unguarded(15) <= ptr_deref_1741_store_0_req_0;
      reqL_unguarded(14) <= ptr_deref_1076_store_0_req_0;
      reqL_unguarded(13) <= ptr_deref_1184_store_0_req_0;
      reqL_unguarded(12) <= ptr_deref_3321_store_0_req_0;
      reqL_unguarded(11) <= ptr_deref_1633_store_0_req_0;
      reqL_unguarded(10) <= ptr_deref_2189_store_0_req_0;
      reqL_unguarded(9) <= ptr_deref_4465_store_0_req_0;
      reqL_unguarded(8) <= ptr_deref_2297_store_0_req_0;
      reqL_unguarded(7) <= ptr_deref_4011_store_0_req_0;
      reqL_unguarded(6) <= ptr_deref_2759_store_0_req_0;
      reqL_unguarded(5) <= ptr_deref_2867_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_3429_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_5029_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_5137_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_3903_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_4573_store_0_req_0;
      ptr_deref_1741_store_0_ack_0 <= ackL_unguarded(15);
      ptr_deref_1076_store_0_ack_0 <= ackL_unguarded(14);
      ptr_deref_1184_store_0_ack_0 <= ackL_unguarded(13);
      ptr_deref_3321_store_0_ack_0 <= ackL_unguarded(12);
      ptr_deref_1633_store_0_ack_0 <= ackL_unguarded(11);
      ptr_deref_2189_store_0_ack_0 <= ackL_unguarded(10);
      ptr_deref_4465_store_0_ack_0 <= ackL_unguarded(9);
      ptr_deref_2297_store_0_ack_0 <= ackL_unguarded(8);
      ptr_deref_4011_store_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_2759_store_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_2867_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_3429_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_5029_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_5137_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_3903_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_4573_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= ptr_deref_1741_store_0_req_1;
      reqR_unguarded(14) <= ptr_deref_1076_store_0_req_1;
      reqR_unguarded(13) <= ptr_deref_1184_store_0_req_1;
      reqR_unguarded(12) <= ptr_deref_3321_store_0_req_1;
      reqR_unguarded(11) <= ptr_deref_1633_store_0_req_1;
      reqR_unguarded(10) <= ptr_deref_2189_store_0_req_1;
      reqR_unguarded(9) <= ptr_deref_4465_store_0_req_1;
      reqR_unguarded(8) <= ptr_deref_2297_store_0_req_1;
      reqR_unguarded(7) <= ptr_deref_4011_store_0_req_1;
      reqR_unguarded(6) <= ptr_deref_2759_store_0_req_1;
      reqR_unguarded(5) <= ptr_deref_2867_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_3429_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_5029_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_5137_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_3903_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_4573_store_0_req_1;
      ptr_deref_1741_store_0_ack_1 <= ackR_unguarded(15);
      ptr_deref_1076_store_0_ack_1 <= ackR_unguarded(14);
      ptr_deref_1184_store_0_ack_1 <= ackR_unguarded(13);
      ptr_deref_3321_store_0_ack_1 <= ackR_unguarded(12);
      ptr_deref_1633_store_0_ack_1 <= ackR_unguarded(11);
      ptr_deref_2189_store_0_ack_1 <= ackR_unguarded(10);
      ptr_deref_4465_store_0_ack_1 <= ackR_unguarded(9);
      ptr_deref_2297_store_0_ack_1 <= ackR_unguarded(8);
      ptr_deref_4011_store_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_2759_store_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_2867_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_3429_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_5029_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_5137_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_3903_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_4573_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      StoreGroup3_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_6: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_7: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_8: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_9: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_10: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_11: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_12: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_13: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_14: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_15: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1741_word_address_0 & ptr_deref_1076_word_address_0 & ptr_deref_1184_word_address_0 & ptr_deref_3321_word_address_0 & ptr_deref_1633_word_address_0 & ptr_deref_2189_word_address_0 & ptr_deref_4465_word_address_0 & ptr_deref_2297_word_address_0 & ptr_deref_4011_word_address_0 & ptr_deref_2759_word_address_0 & ptr_deref_2867_word_address_0 & ptr_deref_3429_word_address_0 & ptr_deref_5029_word_address_0 & ptr_deref_5137_word_address_0 & ptr_deref_3903_word_address_0 & ptr_deref_4573_word_address_0;
      data_in <= ptr_deref_1741_data_0 & ptr_deref_1076_data_0 & ptr_deref_1184_data_0 & ptr_deref_3321_data_0 & ptr_deref_1633_data_0 & ptr_deref_2189_data_0 & ptr_deref_4465_data_0 & ptr_deref_2297_data_0 & ptr_deref_4011_data_0 & ptr_deref_2759_data_0 & ptr_deref_2867_data_0 & ptr_deref_3429_data_0 & ptr_deref_5029_data_0 & ptr_deref_5137_data_0 & ptr_deref_3903_data_0 & ptr_deref_4573_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 16,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared call operator group (0) : call_stmt_5270_call 
    sendOutput_call_group_0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_5270_call_req_0;
      call_stmt_5270_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_5270_call_req_1;
      call_stmt_5270_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_0_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_716_call 
    testConfigure_call_group_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_716_call_req_0;
      call_stmt_716_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_716_call_req_1;
      call_stmt_716_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_1_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_716 <= data_out(15 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          dataL => testConfigure_return_data(15 downto 0),
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    zeropad_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    zeropad_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    zeropad_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(21 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(21 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(21 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(1 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(43 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(9 downto 0);
  -- interface signals to connect to memory space memory_space_3
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(1 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(41 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(7 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(37 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(43 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(9 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(21 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_8
  signal memory_space_8_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_tag : std_logic_vector(21 downto 0);
  signal memory_space_8_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_8_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_8_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(1 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(43 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(9 downto 0);
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(4 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(4 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal testConfigure_out_args   : std_logic_vector(15 downto 0);
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_data: std_logic_vector(15 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module zeropad3D
  component zeropad3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(4 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_data : in   std_logic_vector(15 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D
  signal zeropad3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_start_req : std_logic;
  signal zeropad3D_start_ack : std_logic;
  signal zeropad3D_fin_req   : std_logic;
  signal zeropad3D_fin_ack : std_logic;
  -- aggregate signals for read from pipe zeropad_input_pipe
  signal zeropad_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal zeropad_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal zeropad_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe zeropad_output_pipe
  signal zeropad_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal zeropad_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal zeropad_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(21 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(4 downto 0),
      memory_space_6_lr_req => memory_space_6_lr_req(1 downto 1),
      memory_space_6_lr_ack => memory_space_6_lr_ack(1 downto 1),
      memory_space_6_lr_addr => memory_space_6_lr_addr(13 downto 7),
      memory_space_6_lr_tag => memory_space_6_lr_tag(43 downto 22),
      memory_space_6_lc_req => memory_space_6_lc_req(1 downto 1),
      memory_space_6_lc_ack => memory_space_6_lc_ack(1 downto 1),
      memory_space_6_lc_data => memory_space_6_lc_data(63 downto 32),
      memory_space_6_lc_tag => memory_space_6_lc_tag(9 downto 5),
      zeropad_output_pipe_pipe_write_req => zeropad_output_pipe_pipe_write_req(0 downto 0),
      zeropad_output_pipe_pipe_write_ack => zeropad_output_pipe_pipe_write_ack(0 downto 0),
      zeropad_output_pipe_pipe_write_data => zeropad_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module testConfigure
  testConfigure_out_args <= testConfigure_ret_val_x_x ;
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      return_data =>testConfigure_return_data,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      return_mdata => testConfigure_out_args,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => testConfigure_ret_val_x_x,
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(1 downto 1),
      memory_space_5_lr_ack => memory_space_5_lr_ack(1 downto 1),
      memory_space_5_lr_addr => memory_space_5_lr_addr(13 downto 7),
      memory_space_5_lr_tag => memory_space_5_lr_tag(37 downto 19),
      memory_space_5_lc_req => memory_space_5_lc_req(1 downto 1),
      memory_space_5_lc_ack => memory_space_5_lc_ack(1 downto 1),
      memory_space_5_lc_data => memory_space_5_lc_data(63 downto 32),
      memory_space_5_lc_tag => memory_space_5_lc_tag(3 downto 2),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(20 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(3 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(1 downto 1),
      memory_space_2_sr_ack => memory_space_2_sr_ack(1 downto 1),
      memory_space_2_sr_addr => memory_space_2_sr_addr(1 downto 1),
      memory_space_2_sr_data => memory_space_2_sr_data(15 downto 8),
      memory_space_2_sr_tag => memory_space_2_sr_tag(43 downto 22),
      memory_space_2_sc_req => memory_space_2_sc_req(1 downto 1),
      memory_space_2_sc_ack => memory_space_2_sc_ack(1 downto 1),
      memory_space_2_sc_tag => memory_space_2_sc_tag(9 downto 5),
      memory_space_4_sr_req => memory_space_4_sr_req(1 downto 1),
      memory_space_4_sr_ack => memory_space_4_sr_ack(1 downto 1),
      memory_space_4_sr_addr => memory_space_4_sr_addr(1 downto 1),
      memory_space_4_sr_data => memory_space_4_sr_data(15 downto 8),
      memory_space_4_sr_tag => memory_space_4_sr_tag(41 downto 21),
      memory_space_4_sc_req => memory_space_4_sc_req(1 downto 1),
      memory_space_4_sc_ack => memory_space_4_sc_ack(1 downto 1),
      memory_space_4_sc_tag => memory_space_4_sc_tag(7 downto 4),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(6 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(31 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(18 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(1 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(6 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(31 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(21 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(4 downto 0),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(7 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(20 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(3 downto 0),
      memory_space_8_sr_req => memory_space_8_sr_req(1 downto 1),
      memory_space_8_sr_ack => memory_space_8_sr_ack(1 downto 1),
      memory_space_8_sr_addr => memory_space_8_sr_addr(1 downto 1),
      memory_space_8_sr_data => memory_space_8_sr_data(15 downto 8),
      memory_space_8_sr_tag => memory_space_8_sr_tag(43 downto 22),
      memory_space_8_sc_req => memory_space_8_sc_req(1 downto 1),
      memory_space_8_sc_ack => memory_space_8_sc_ack(1 downto 1),
      memory_space_8_sc_tag => memory_space_8_sc_tag(9 downto 5),
      zeropad_input_pipe_pipe_read_req => zeropad_input_pipe_pipe_read_req(0 downto 0),
      zeropad_input_pipe_pipe_read_ack => zeropad_input_pipe_pipe_read_ack(0 downto 0),
      zeropad_input_pipe_pipe_read_data => zeropad_input_pipe_pipe_read_data(7 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  -- module zeropad3D
  zeropad3D_instance:zeropad3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_start_req,
      start_ack => zeropad3D_start_ack,
      fin_req => zeropad3D_fin_req,
      fin_ack => zeropad3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(20 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(21 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(7 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(4 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(0 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(20 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(7 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(3 downto 0),
      memory_space_5_lr_req => memory_space_5_lr_req(0 downto 0),
      memory_space_5_lr_ack => memory_space_5_lr_ack(0 downto 0),
      memory_space_5_lr_addr => memory_space_5_lr_addr(6 downto 0),
      memory_space_5_lr_tag => memory_space_5_lr_tag(18 downto 0),
      memory_space_5_lc_req => memory_space_5_lc_req(0 downto 0),
      memory_space_5_lc_ack => memory_space_5_lc_ack(0 downto 0),
      memory_space_5_lc_data => memory_space_5_lc_data(31 downto 0),
      memory_space_5_lc_tag => memory_space_5_lc_tag(1 downto 0),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(6 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(21 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(31 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(4 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(20 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(7 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(3 downto 0),
      memory_space_8_lr_req => memory_space_8_lr_req(0 downto 0),
      memory_space_8_lr_ack => memory_space_8_lr_ack(0 downto 0),
      memory_space_8_lr_addr => memory_space_8_lr_addr(0 downto 0),
      memory_space_8_lr_tag => memory_space_8_lr_tag(21 downto 0),
      memory_space_8_lc_req => memory_space_8_lc_req(0 downto 0),
      memory_space_8_lc_ack => memory_space_8_lc_ack(0 downto 0),
      memory_space_8_lc_data => memory_space_8_lc_data(7 downto 0),
      memory_space_8_lc_tag => memory_space_8_lc_tag(4 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(21 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(4 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(7 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(21 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(4 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(0 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(7 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(20 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(3 downto 0),
      memory_space_8_sr_req => memory_space_8_sr_req(0 downto 0),
      memory_space_8_sr_ack => memory_space_8_sr_ack(0 downto 0),
      memory_space_8_sr_addr => memory_space_8_sr_addr(0 downto 0),
      memory_space_8_sr_data => memory_space_8_sr_data(7 downto 0),
      memory_space_8_sr_tag => memory_space_8_sr_tag(21 downto 0),
      memory_space_8_sc_req => memory_space_8_sc_req(0 downto 0),
      memory_space_8_sc_ack => memory_space_8_sc_ack(0 downto 0),
      memory_space_8_sc_tag => memory_space_8_sc_tag(4 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_data => testConfigure_return_data(15 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      tag_in => zeropad3D_tag_in,
      tag_out => zeropad3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_tag_in <= (others => '0');
  zeropad3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_start_req, start_ack => zeropad3D_start_ack,  fin_req => zeropad3D_fin_req,  fin_ack => zeropad3D_fin_ack);
  zeropad_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_input_pipe_pipe_read_req,
      read_ack => zeropad_input_pipe_pipe_read_ack,
      read_data => zeropad_input_pipe_pipe_read_data,
      write_req => zeropad_input_pipe_pipe_write_req,
      write_ack => zeropad_input_pipe_pipe_write_ack,
      write_data => zeropad_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_output_pipe_pipe_read_req,
      read_ack => zeropad_output_pipe_pipe_read_ack,
      read_data => zeropad_output_pipe_pipe_read_data,
      write_req => zeropad_output_pipe_pipe_write_req,
      write_ack => zeropad_output_pipe_pipe_write_ack,
      write_data => zeropad_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 2,
      addr_width => 1,
      data_width => 8,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 1,
      num_stores => 2,
      addr_width => 1,
      data_width => 8,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_loads => 2,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 2,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_8: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_8",
      num_loads => 1,
      num_stores => 2,
      addr_width => 1,
      data_width => 8,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_8_lr_addr,
      lr_req_in => memory_space_8_lr_req,
      lr_ack_out => memory_space_8_lr_ack,
      lr_tag_in => memory_space_8_lr_tag,
      lc_req_in => memory_space_8_lc_req,
      lc_ack_out => memory_space_8_lc_ack,
      lc_data_out => memory_space_8_lc_data,
      lc_tag_out => memory_space_8_lc_tag,
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
