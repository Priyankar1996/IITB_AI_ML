-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    num_cont : in  std_logic_vector(15 downto 0);
    row1 : in  std_logic_vector(15 downto 0);
    col1 : in  std_logic_vector(15 downto 0);
    rk1 : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 96)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal num_cont_buffer :  std_logic_vector(15 downto 0);
  signal num_cont_update_enable: Boolean;
  signal row1_buffer :  std_logic_vector(15 downto 0);
  signal row1_update_enable: Boolean;
  signal col1_buffer :  std_logic_vector(15 downto 0);
  signal col1_update_enable: Boolean;
  signal rk1_buffer :  std_logic_vector(15 downto 0);
  signal rk1_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_43_branch_req_0 : boolean;
  signal phi_stmt_45_ack_0 : boolean;
  signal phi_stmt_45_req_0 : boolean;
  signal phi_stmt_45_req_1 : boolean;
  signal n_address_279_47_buf_req_0 : boolean;
  signal n_address_279_47_buf_ack_0 : boolean;
  signal n_address_279_47_buf_req_1 : boolean;
  signal n_address_279_47_buf_ack_1 : boolean;
  signal phi_stmt_50_req_0 : boolean;
  signal phi_stmt_50_req_1 : boolean;
  signal phi_stmt_50_ack_0 : boolean;
  signal n_word_start_268_52_buf_req_0 : boolean;
  signal n_word_start_268_52_buf_ack_0 : boolean;
  signal n_word_start_268_52_buf_req_1 : boolean;
  signal n_word_start_268_52_buf_ack_1 : boolean;
  signal n_winr_208_69_buf_req_0 : boolean;
  signal n_winr_208_69_buf_ack_0 : boolean;
  signal phi_stmt_56_req_1 : boolean;
  signal phi_stmt_56_req_0 : boolean;
  signal phi_stmt_56_ack_0 : boolean;
  signal nl_start_34_58_buf_req_0 : boolean;
  signal nl_start_34_58_buf_ack_0 : boolean;
  signal nl_start_34_58_buf_req_1 : boolean;
  signal nl_start_34_58_buf_ack_1 : boolean;
  signal n_left_287_59_buf_req_0 : boolean;
  signal n_left_287_59_buf_ack_0 : boolean;
  signal n_left_287_59_buf_req_1 : boolean;
  signal n_left_287_59_buf_ack_1 : boolean;
  signal phi_stmt_60_req_0 : boolean;
  signal phi_stmt_60_req_1 : boolean;
  signal phi_stmt_60_ack_0 : boolean;
  signal n_blk_307_62_buf_req_0 : boolean;
  signal n_blk_307_62_buf_ack_0 : boolean;
  signal n_blk_307_62_buf_req_1 : boolean;
  signal n_blk_307_62_buf_ack_1 : boolean;
  signal type_cast_64_inst_req_0 : boolean;
  signal type_cast_64_inst_ack_0 : boolean;
  signal type_cast_64_inst_req_1 : boolean;
  signal type_cast_64_inst_ack_1 : boolean;
  signal phi_stmt_65_req_1 : boolean;
  signal phi_stmt_65_req_0 : boolean;
  signal phi_stmt_65_ack_0 : boolean;
  signal WPIPE_input_pipe1_166_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_166_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_166_inst_ack_1 : boolean;
  signal W_c3_163_delayed_14_0_169_inst_req_0 : boolean;
  signal W_c3_163_delayed_14_0_169_inst_ack_0 : boolean;
  signal W_c3_163_delayed_14_0_169_inst_req_1 : boolean;
  signal W_c3_163_delayed_14_0_169_inst_ack_1 : boolean;
  signal n_winr_208_69_buf_req_1 : boolean;
  signal n_winr_208_69_buf_ack_1 : boolean;
  signal phi_stmt_70_req_1 : boolean;
  signal phi_stmt_70_req_0 : boolean;
  signal phi_stmt_70_ack_0 : boolean;
  signal n_col_221_74_buf_req_0 : boolean;
  signal n_col_221_74_buf_ack_0 : boolean;
  signal n_col_221_74_buf_req_1 : boolean;
  signal n_col_221_74_buf_ack_1 : boolean;
  signal phi_stmt_75_req_0 : boolean;
  signal phi_stmt_75_req_1 : boolean;
  signal phi_stmt_75_ack_0 : boolean;
  signal n_row_233_77_buf_req_0 : boolean;
  signal n_row_233_77_buf_ack_0 : boolean;
  signal n_row_233_77_buf_req_1 : boolean;
  signal n_row_233_77_buf_ack_1 : boolean;
  signal array_obj_ref_132_index_offset_req_0 : boolean;
  signal array_obj_ref_132_index_offset_ack_0 : boolean;
  signal array_obj_ref_132_index_offset_req_1 : boolean;
  signal array_obj_ref_132_index_offset_ack_1 : boolean;
  signal addr_of_133_final_reg_req_0 : boolean;
  signal addr_of_133_final_reg_ack_0 : boolean;
  signal addr_of_133_final_reg_req_1 : boolean;
  signal addr_of_133_final_reg_ack_1 : boolean;
  signal ptr_deref_137_load_0_req_0 : boolean;
  signal ptr_deref_137_load_0_ack_0 : boolean;
  signal ptr_deref_137_load_0_req_1 : boolean;
  signal ptr_deref_137_load_0_ack_1 : boolean;
  signal slice_141_inst_req_0 : boolean;
  signal slice_141_inst_ack_0 : boolean;
  signal slice_141_inst_req_1 : boolean;
  signal slice_141_inst_ack_1 : boolean;
  signal slice_145_inst_req_0 : boolean;
  signal slice_145_inst_ack_0 : boolean;
  signal slice_145_inst_req_1 : boolean;
  signal slice_145_inst_ack_1 : boolean;
  signal slice_149_inst_req_0 : boolean;
  signal slice_149_inst_ack_0 : boolean;
  signal slice_149_inst_req_1 : boolean;
  signal slice_149_inst_ack_1 : boolean;
  signal slice_153_inst_req_0 : boolean;
  signal slice_153_inst_ack_0 : boolean;
  signal slice_153_inst_req_1 : boolean;
  signal slice_153_inst_ack_1 : boolean;
  signal W_c1_155_delayed_14_0_155_inst_req_0 : boolean;
  signal W_c1_155_delayed_14_0_155_inst_ack_0 : boolean;
  signal W_c1_155_delayed_14_0_155_inst_req_1 : boolean;
  signal W_c1_155_delayed_14_0_155_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_159_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_159_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_159_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_159_inst_ack_1 : boolean;
  signal W_c2_159_delayed_14_0_162_inst_req_0 : boolean;
  signal W_c2_159_delayed_14_0_162_inst_ack_0 : boolean;
  signal W_c2_159_delayed_14_0_162_inst_req_1 : boolean;
  signal W_c2_159_delayed_14_0_162_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_166_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_173_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_173_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_173_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_173_inst_ack_1 : boolean;
  signal W_c4_167_delayed_14_0_176_inst_req_0 : boolean;
  signal W_c4_167_delayed_14_0_176_inst_ack_0 : boolean;
  signal W_c4_167_delayed_14_0_176_inst_req_1 : boolean;
  signal W_c4_167_delayed_14_0_176_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_180_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_180_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_180_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_180_inst_ack_1 : boolean;
  signal do_while_stmt_43_branch_ack_0 : boolean;
  signal do_while_stmt_43_branch_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 96) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= num_cont;
  num_cont_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= row1;
  row1_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= col1;
  col1_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(63 downto 48) <= rk1;
  rk1_buffer <= in_buffer_data_out(63 downto 48);
  in_buffer_data_in(79 downto 64) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(95 downto 80) <= ct;
  ct_buffer <= in_buffer_data_out(95 downto 80);
  in_buffer_data_in(tag_length + 95 downto 96) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 95 downto 96);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,access_T_CP_0_start,"access_T cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,access_T_CP_0_symbol, "access_T cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(207 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_31_to_assign_stmt_42__exit__
      -- CP-element group 0: 	 branch_block_stmt_25/do_while_stmt_43__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_25/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/branch_block_stmt_25__entry__
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_31_to_assign_stmt_42__entry__
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_31_to_assign_stmt_42/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_31_to_assign_stmt_42/$exit
      -- 
    -- logger for CP element group access_T_CP_0_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	207 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_25/$exit
      -- CP-element group 1: 	 branch_block_stmt_25/branch_block_stmt_25__exit__
      -- CP-element group 1: 	 branch_block_stmt_25/do_while_stmt_43__exit__
      -- 
    -- logger for CP element group access_T_CP_0_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(207);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_25/do_while_stmt_43/$entry
      -- CP-element group 2: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43__entry__
      -- 
    -- logger for CP element group access_T_CP_0_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(2) <= access_T_CP_0_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	207 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43__exit__
      -- 
    -- logger for CP element group access_T_CP_0_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_25/do_while_stmt_43/loop_back
      -- 
    -- logger for CP element group access_T_CP_0_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	205 
    -- CP-element group 5: 	206 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_25/do_while_stmt_43/condition_done
      -- CP-element group 5: 	 branch_block_stmt_25/do_while_stmt_43/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_25/do_while_stmt_43/loop_taken/$entry
      -- 
    -- logger for CP element group access_T_CP_0_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(5) <= access_T_CP_0_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	204 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_25/do_while_stmt_43/loop_body_done
      -- 
    -- logger for CP element group access_T_CP_0_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(6) <= access_T_CP_0_elements(204);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	38 
    -- CP-element group 7: 	76 
    -- CP-element group 7: 	97 
    -- CP-element group 7: 	116 
    -- CP-element group 7: 	135 
    -- CP-element group 7: 	57 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group access_T_CP_0_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(7) <= access_T_CP_0_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	40 
    -- CP-element group 8: 	78 
    -- CP-element group 8: 	99 
    -- CP-element group 8: 	118 
    -- CP-element group 8: 	137 
    -- CP-element group 8: 	59 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group access_T_CP_0_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(8) <= access_T_CP_0_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	70 
    -- CP-element group 9: 	71 
    -- CP-element group 9: 	91 
    -- CP-element group 9: 	92 
    -- CP-element group 9: 	110 
    -- CP-element group 9: 	111 
    -- CP-element group 9: 	129 
    -- CP-element group 9: 	130 
    -- CP-element group 9: 	149 
    -- CP-element group 9: 	150 
    -- CP-element group 9: 	203 
    -- CP-element group 9: 	51 
    -- CP-element group 9: 	52 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/loop_body_start
      -- 
    -- logger for CP element group access_T_CP_0_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	203 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/condition_evaluated
      -- 
    -- logger for CP element group access_T_CP_0_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:do_while_stmt_43_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(10), ack => do_while_stmt_43_branch_req_0); -- 
    access_T_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(14) & access_T_CP_0_elements(203);
      gj_access_T_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	70 
    -- CP-element group 11: 	91 
    -- CP-element group 11: 	110 
    -- CP-element group 11: 	129 
    -- CP-element group 11: 	51 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	72 
    -- CP-element group 11: 	93 
    -- CP-element group 11: 	112 
    -- CP-element group 11: 	131 
    -- CP-element group 11: 	53 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_sample_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= access_T_CP_0_elements(15) & access_T_CP_0_elements(32) & access_T_CP_0_elements(70) & access_T_CP_0_elements(91) & access_T_CP_0_elements(110) & access_T_CP_0_elements(129) & access_T_CP_0_elements(51) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	73 
    -- CP-element group 12: 	94 
    -- CP-element group 12: 	113 
    -- CP-element group 12: 	132 
    -- CP-element group 12: 	54 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	204 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	32 
    -- CP-element group 12: 	70 
    -- CP-element group 12: 	91 
    -- CP-element group 12: 	110 
    -- CP-element group 12: 	129 
    -- CP-element group 12: 	51 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_sample_completed_
      -- 
    -- logger for CP element group access_T_CP_0_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(17) & access_T_CP_0_elements(35) & access_T_CP_0_elements(73) & access_T_CP_0_elements(94) & access_T_CP_0_elements(113) & access_T_CP_0_elements(132) & access_T_CP_0_elements(54);
      gj_access_T_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	33 
    -- CP-element group 13: 	71 
    -- CP-element group 13: 	92 
    -- CP-element group 13: 	111 
    -- CP-element group 13: 	130 
    -- CP-element group 13: 	52 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	74 
    -- CP-element group 13: 	95 
    -- CP-element group 13: 	114 
    -- CP-element group 13: 	133 
    -- CP-element group 13: 	55 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_update_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(16) & access_T_CP_0_elements(33) & access_T_CP_0_elements(71) & access_T_CP_0_elements(92) & access_T_CP_0_elements(111) & access_T_CP_0_elements(130) & access_T_CP_0_elements(52);
      gj_access_T_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	96 
    -- CP-element group 14: 	115 
    -- CP-element group 14: 	134 
    -- CP-element group 14: 	56 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(18) & access_T_CP_0_elements(37) & access_T_CP_0_elements(75) & access_T_CP_0_elements(96) & access_T_CP_0_elements(115) & access_T_CP_0_elements(134) & access_T_CP_0_elements(56);
      gj_access_T_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_sample_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	151 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_update_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(151);
      gj_access_T_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_sample_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	151 
    -- CP-element group 18:  members (15) 
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_index_resized_1
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_index_scaled_1
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_index_computed_1
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_index_resize_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_index_resize_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_index_resize_1/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_index_resize_1/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_index_scale_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_index_scale_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_index_scale_1/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_index_scale_1/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_final_index_sum_regn_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_final_index_sum_regn_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:array_obj_ref_132_index_offset_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(18), ack => array_obj_ref_132_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_loopback_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(19) <= access_T_CP_0_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_loopback_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_45_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_45_loopback_sample_req_44_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_45_loopback_sample_req_44_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(20), ack => phi_stmt_45_req_0); -- 
    -- Element group access_T_CP_0_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_entry_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(21) <= access_T_CP_0_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_entry_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_45_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_45_entry_sample_req_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_45_entry_sample_req_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(22), ack => phi_stmt_45_req_1); -- 
    -- Element group access_T_CP_0_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_45_phi_mux_ack_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_45_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_45_phi_mux_ack_50_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_45_ack_0, ack => access_T_CP_0_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_address_279_47_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_63_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_63_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(24), ack => n_address_279_47_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_update_start_
      -- CP-element group 25: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_address_279_47_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_68_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_68_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(25), ack => n_address_279_47_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_Sample/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_address_279_47_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_64_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_279_47_buf_ack_0, ack => access_T_CP_0_elements(26)); -- 
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_address_47_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_address_279_47_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_69_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_279_47_buf_ack_1, ack => access_T_CP_0_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_49_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_49_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_49_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_49_sample_completed_
      -- 
    -- logger for CP element group access_T_CP_0_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(28) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_49_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_49_update_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(29) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_49_update_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(30) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(30) <= access_T_CP_0_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_49_update_completed_
      -- 
    -- logger for CP element group access_T_CP_0_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(31) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(29), ack => access_T_CP_0_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	12 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_sample_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(32) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	177 
    -- CP-element group 33: 	184 
    -- CP-element group 33: 	191 
    -- CP-element group 33: 	198 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_update_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(33) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(177) & access_T_CP_0_elements(184) & access_T_CP_0_elements(191) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_sample_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(34) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(34) <= access_T_CP_0_elements(11);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_sample_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(35) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_update_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(36) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(36) <= access_T_CP_0_elements(13);
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: 	175 
    -- CP-element group 37: 	182 
    -- CP-element group 37: 	189 
    -- CP-element group 37: 	196 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_update_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(37) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_loopback_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(38) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_loopback_sample_req
      -- CP-element group 39: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_loopback_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_50_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_50_loopback_sample_req_88_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_50_loopback_sample_req_88_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(39), ack => phi_stmt_50_req_0); -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_entry_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(40) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(40) <= access_T_CP_0_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_entry_sample_req
      -- CP-element group 41: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_entry_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_50_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_50_entry_sample_req_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_50_entry_sample_req_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(41), ack => phi_stmt_50_req_1); -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_phi_mux_ack
      -- CP-element group 42: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_50_phi_mux_ack_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_50_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_50_phi_mux_ack_94_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_50_ack_0, ack => access_T_CP_0_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_sample_start__ps
      -- CP-element group 43: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_word_start_268_52_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(43), ack => n_word_start_268_52_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_update_start__ps
      -- CP-element group 44: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_update_start_
      -- CP-element group 44: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_word_start_268_52_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(44), ack => n_word_start_268_52_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_Sample/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_word_start_268_52_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_268_52_buf_ack_0, ack => access_T_CP_0_elements(45)); -- 
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_update_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_word_start_52_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_word_start_268_52_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_268_52_buf_ack_1, ack => access_T_CP_0_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_55_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_55_sample_completed__ps
      -- CP-element group 47: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_55_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_55_sample_completed_
      -- 
    -- logger for CP element group access_T_CP_0_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(47) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_55_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_55_update_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(48) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_55_update_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(49) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(49) <= access_T_CP_0_elements(50);
    -- CP-element group 50:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	49 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_55_update_completed_
      -- 
    -- logger for CP element group access_T_CP_0_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(50) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(50) is a control-delay.
    cp_element_50_delay: control_delay_element  generic map(name => " 50_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(48), ack => access_T_CP_0_elements(50), clk => clk, reset =>reset);
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	9 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	12 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	11 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_sample_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(51) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	9 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	56 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	13 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_update_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(52) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(56);
      gj_access_T_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_sample_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(53) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(53) <= access_T_CP_0_elements(11);
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	12 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_sample_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(54) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_update_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(55) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(55) <= access_T_CP_0_elements(13);
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	14 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	52 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_update_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(56) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	7 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_loopback_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(57) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(57) <= access_T_CP_0_elements(7);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_loopback_sample_req
      -- CP-element group 58: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_loopback_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_56_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_56_loopback_sample_req_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_56_loopback_sample_req_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(58), ack => phi_stmt_56_req_1); -- 
    -- Element group access_T_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	8 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_entry_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(59) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(59) <= access_T_CP_0_elements(8);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_entry_sample_req
      -- CP-element group 60: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_entry_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_56_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_56_entry_sample_req_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_56_entry_sample_req_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(60), ack => phi_stmt_56_req_0); -- 
    -- Element group access_T_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_phi_mux_ack
      -- CP-element group 61: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_56_phi_mux_ack_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_56_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_56_phi_mux_ack_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_56_ack_0, ack => access_T_CP_0_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_sample_start__ps
      -- CP-element group 62: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:nl_start_34_58_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(62), ack => nl_start_34_58_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_update_start__ps
      -- CP-element group 63: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_update_start_
      -- CP-element group 63: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:nl_start_34_58_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(63), ack => nl_start_34_58_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_sample_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_Sample/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:nl_start_34_58_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_34_58_buf_ack_0, ack => access_T_CP_0_elements(64)); -- 
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_update_completed__ps
      -- CP-element group 65: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_nl_start_58_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:nl_start_34_58_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_34_58_buf_ack_1, ack => access_T_CP_0_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_left_287_59_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(66), ack => n_left_287_59_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_update_start_
      -- CP-element group 67: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_left_287_59_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(67), ack => n_left_287_59_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_Sample/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_left_287_59_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_287_59_buf_ack_0, ack => access_T_CP_0_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_left_59_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_left_287_59_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_287_59_buf_ack_1, ack => access_T_CP_0_elements(69)); -- 
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	9 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	12 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	11 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_sample_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(70) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	9 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	184 
    -- CP-element group 71: 	191 
    -- CP-element group 71: 	198 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	13 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_update_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(71) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(184) & access_T_CP_0_elements(191) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_sample_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(72) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(72) <= access_T_CP_0_elements(11);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	12 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_sample_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(73) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	13 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_update_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(74) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(74) <= access_T_CP_0_elements(13);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: 	182 
    -- CP-element group 75: 	189 
    -- CP-element group 75: 	196 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_update_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(75) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	7 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_loopback_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(76) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(76) <= access_T_CP_0_elements(7);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_loopback_sample_req
      -- CP-element group 77: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_loopback_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_60_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_60_loopback_sample_req_186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_60_loopback_sample_req_186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(77), ack => phi_stmt_60_req_0); -- 
    -- Element group access_T_CP_0_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	8 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_entry_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(78) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(78) <= access_T_CP_0_elements(8);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_entry_sample_req
      -- CP-element group 79: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_entry_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_60_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_60_entry_sample_req_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_60_entry_sample_req_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(79), ack => phi_stmt_60_req_1); -- 
    -- Element group access_T_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_phi_mux_ack
      -- CP-element group 80: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_60_phi_mux_ack_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_60_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_60_phi_mux_ack_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_60_ack_0, ack => access_T_CP_0_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_sample_start__ps
      -- CP-element group 81: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(81) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_blk_307_62_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(81), ack => n_blk_307_62_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_update_start__ps
      -- CP-element group 82: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_update_start_
      -- CP-element group 82: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_blk_307_62_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(82), ack => n_blk_307_62_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_sample_completed__ps
      -- CP-element group 83: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_Sample/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(83) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_blk_307_62_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_307_62_buf_ack_0, ack => access_T_CP_0_elements(83)); -- 
    -- CP-element group 84:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_update_completed__ps
      -- CP-element group 84: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_blk_62_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(84) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_blk_307_62_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_307_62_buf_ack_1, ack => access_T_CP_0_elements(84)); -- 
    -- CP-element group 85:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_sample_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(85) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_update_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(86) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	89 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_Sample/rr
      -- 
    -- logger for CP element group access_T_CP_0_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(87) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:type_cast_64_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(87), ack => type_cast_64_inst_req_0); -- 
    access_T_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(85) & access_T_CP_0_elements(89);
      gj_access_T_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_update_start_
      -- CP-element group 88: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_Update/cr
      -- 
    -- logger for CP element group access_T_CP_0_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:type_cast_64_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(88), ack => type_cast_64_inst_req_1); -- 
    access_T_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(86) & access_T_CP_0_elements(90);
      gj_access_T_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	87 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_Sample/ra
      -- 
    -- logger for CP element group access_T_CP_0_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:type_cast_64_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_0, ack => access_T_CP_0_elements(89)); -- 
    -- CP-element group 90:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_update_completed__ps
      -- CP-element group 90: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_64_Update/ca
      -- 
    -- logger for CP element group access_T_CP_0_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(90) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:type_cast_64_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_1, ack => access_T_CP_0_elements(90)); -- 
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	9 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	12 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	11 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_sample_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(91) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	9 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	96 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	13 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_update_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(92) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(96);
      gj_access_T_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	11 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_sample_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(93) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(93) <= access_T_CP_0_elements(11);
    -- CP-element group 94:  join  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	12 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_sample_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(94) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(94) is bound as output of CP function.
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	13 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_update_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(95) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(95) <= access_T_CP_0_elements(13);
    -- CP-element group 96:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	14 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	92 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_update_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(96) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	7 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_loopback_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(97) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(97) <= access_T_CP_0_elements(7);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_loopback_sample_req
      -- CP-element group 98: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_loopback_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_65_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_65_loopback_sample_req_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_65_loopback_sample_req_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(98), ack => phi_stmt_65_req_1); -- 
    -- Element group access_T_CP_0_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	8 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_entry_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(99) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(99) <= access_T_CP_0_elements(8);
    -- CP-element group 100:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_entry_sample_req
      -- CP-element group 100: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_entry_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(100) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_65_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_65_entry_sample_req_243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_65_entry_sample_req_243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(100), ack => phi_stmt_65_req_0); -- 
    -- Element group access_T_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_phi_mux_ack
      -- CP-element group 101: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_65_phi_mux_ack_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(101) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_65_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_65_phi_mux_ack_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_65_ack_0, ack => access_T_CP_0_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_68_sample_start__ps
      -- CP-element group 102: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_68_sample_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_68_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_68_sample_completed_
      -- 
    -- logger for CP element group access_T_CP_0_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(102) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_68_update_start__ps
      -- CP-element group 103: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_68_update_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(103) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(103) is bound as output of CP function.
    -- CP-element group 104:  join  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_68_update_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(104) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(104) <= access_T_CP_0_elements(105);
    -- CP-element group 105:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	104 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_68_update_completed_
      -- 
    -- logger for CP element group access_T_CP_0_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(105) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(103), ack => access_T_CP_0_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_sample_start__ps
      -- CP-element group 106: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(106) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_winr_208_69_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(106), ack => n_winr_208_69_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_update_start__ps
      -- CP-element group 107: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_update_start_
      -- CP-element group 107: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(107)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(107)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(107) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_winr_208_69_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(107), ack => n_winr_208_69_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_Sample/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(108)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(108)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(108) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_winr_208_69_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_208_69_buf_ack_0, ack => access_T_CP_0_elements(108)); -- 
    -- CP-element group 109:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_update_completed__ps
      -- CP-element group 109: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_winr_69_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(109)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(109)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(109) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_winr_208_69_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_208_69_buf_ack_1, ack => access_T_CP_0_elements(109)); -- 
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	9 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	12 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	11 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_sample_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(110)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(110)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(110) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	9 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	115 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	13 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_update_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(111)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(111)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(111) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(115);
      gj_access_T_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	11 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_sample_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(112)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(112)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(112) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(112) <= access_T_CP_0_elements(11);
    -- CP-element group 113:  join  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	12 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_sample_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(113)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(113)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(113) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(113) is bound as output of CP function.
    -- CP-element group 114:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	13 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_update_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(114)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(114)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(114) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(114) <= access_T_CP_0_elements(13);
    -- CP-element group 115:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	14 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	111 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_update_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(115)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(115)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(115) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(115) is bound as output of CP function.
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	7 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_loopback_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(116)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(116)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(116) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(116) <= access_T_CP_0_elements(7);
    -- CP-element group 117:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_loopback_sample_req
      -- CP-element group 117: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_loopback_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(117)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(117)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(117) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_70_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_70_loopback_sample_req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_70_loopback_sample_req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(117), ack => phi_stmt_70_req_1); -- 
    -- Element group access_T_CP_0_elements(117) is bound as output of CP function.
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	8 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_entry_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(118)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(118)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(118) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(118) <= access_T_CP_0_elements(8);
    -- CP-element group 119:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_entry_sample_req
      -- CP-element group 119: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_entry_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(119)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(119)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(119) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_70_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_70_entry_sample_req_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_70_entry_sample_req_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(119), ack => phi_stmt_70_req_0); -- 
    -- Element group access_T_CP_0_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_phi_mux_ack
      -- CP-element group 120: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_70_phi_mux_ack_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(120)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(120)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(120) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_70_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_70_phi_mux_ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_70_ack_0, ack => access_T_CP_0_elements(120)); -- 
    -- CP-element group 121:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_73_sample_start__ps
      -- CP-element group 121: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_73_sample_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_73_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_73_sample_completed_
      -- 
    -- logger for CP element group access_T_CP_0_elements(121)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(121)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(121) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(121) is bound as output of CP function.
    -- CP-element group 122:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_73_update_start__ps
      -- CP-element group 122: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_73_update_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(122)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(122)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(122) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(122) is bound as output of CP function.
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_73_update_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(123)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(123)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(123) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(123) <= access_T_CP_0_elements(124);
    -- CP-element group 124:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	123 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_73_update_completed_
      -- 
    -- logger for CP element group access_T_CP_0_elements(124)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(124)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(124) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(124) is a control-delay.
    cp_element_124_delay: control_delay_element  generic map(name => " 124_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(122), ack => access_T_CP_0_elements(124), clk => clk, reset =>reset);
    -- CP-element group 125:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_sample_start__ps
      -- CP-element group 125: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(125)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(125)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(125) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_col_221_74_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(125), ack => n_col_221_74_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_update_start__ps
      -- CP-element group 126: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_update_start_
      -- CP-element group 126: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(126)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(126)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(126) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_col_221_74_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(126), ack => n_col_221_74_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(126) is bound as output of CP function.
    -- CP-element group 127:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_Sample/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(127)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(127)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(127) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_col_221_74_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_221_74_buf_ack_0, ack => access_T_CP_0_elements(127)); -- 
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (4) 
      -- CP-element group 128: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_update_completed__ps
      -- CP-element group 128: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_col_74_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(128)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(128)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(128) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_col_221_74_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_221_74_buf_ack_1, ack => access_T_CP_0_elements(128)); -- 
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	9 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	12 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	11 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_sample_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(129)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(129)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(129) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	9 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	134 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	13 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_update_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(130)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(130)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(130) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(134);
      gj_access_T_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	11 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_sample_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(131)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(131)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(131) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(131) <= access_T_CP_0_elements(11);
    -- CP-element group 132:  join  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	12 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_sample_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(132)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(132)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(132) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(132) is bound as output of CP function.
    -- CP-element group 133:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	13 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_update_start__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(133)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(133)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(133) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(133) <= access_T_CP_0_elements(13);
    -- CP-element group 134:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	14 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	130 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_update_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(134)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(134)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(134) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(134) is bound as output of CP function.
    -- CP-element group 135:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	7 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_loopback_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(135)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(135)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(135) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(135) <= access_T_CP_0_elements(7);
    -- CP-element group 136:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_loopback_sample_req
      -- CP-element group 136: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_loopback_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(136)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(136)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(136) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_75_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_75_loopback_sample_req_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_75_loopback_sample_req_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(136), ack => phi_stmt_75_req_0); -- 
    -- Element group access_T_CP_0_elements(136) is bound as output of CP function.
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	8 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_entry_trigger
      -- 
    -- logger for CP element group access_T_CP_0_elements(137)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(137)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(137) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(137) <= access_T_CP_0_elements(8);
    -- CP-element group 138:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_entry_sample_req
      -- CP-element group 138: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_entry_sample_req_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(138)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(138)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(138) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_75_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_75_entry_sample_req_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_75_entry_sample_req_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(138), ack => phi_stmt_75_req_1); -- 
    -- Element group access_T_CP_0_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (2) 
      -- CP-element group 139: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_phi_mux_ack
      -- CP-element group 139: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/phi_stmt_75_phi_mux_ack_ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(139)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(139)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(139) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:phi_stmt_75_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_75_phi_mux_ack_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_75_ack_0, ack => access_T_CP_0_elements(139)); -- 
    -- CP-element group 140:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_sample_start__ps
      -- CP-element group 140: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(140)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(140)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(140) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_row_233_77_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(140), ack => n_row_233_77_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(140) is bound as output of CP function.
    -- CP-element group 141:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (4) 
      -- CP-element group 141: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_update_start__ps
      -- CP-element group 141: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_update_start_
      -- CP-element group 141: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(141)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(141)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(141) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_row_233_77_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(141), ack => n_row_233_77_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(141) is bound as output of CP function.
    -- CP-element group 142:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (4) 
      -- CP-element group 142: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_sample_completed__ps
      -- CP-element group 142: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_Sample/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(142)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(142)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(142) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_row_233_77_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_233_77_buf_ack_0, ack => access_T_CP_0_elements(142)); -- 
    -- CP-element group 143:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (4) 
      -- CP-element group 143: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_update_completed__ps
      -- CP-element group 143: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/R_n_row_77_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(143)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(143)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(143) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:n_row_233_77_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_233_77_buf_ack_1, ack => access_T_CP_0_elements(143)); -- 
    -- CP-element group 144:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_79_sample_start__ps
      -- CP-element group 144: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_79_sample_completed__ps
      -- CP-element group 144: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_79_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_79_sample_completed_
      -- 
    -- logger for CP element group access_T_CP_0_elements(144)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(144)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(144) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_79_update_start__ps
      -- CP-element group 145: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_79_update_start_
      -- 
    -- logger for CP element group access_T_CP_0_elements(145)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(145)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(145) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(145) is bound as output of CP function.
    -- CP-element group 146:  join  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (1) 
      -- CP-element group 146: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_79_update_completed__ps
      -- 
    -- logger for CP element group access_T_CP_0_elements(146)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(146)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(146) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(146) <= access_T_CP_0_elements(147);
    -- CP-element group 147:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	146 
    -- CP-element group 147:  members (1) 
      -- CP-element group 147: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/type_cast_79_update_completed_
      -- 
    -- logger for CP element group access_T_CP_0_elements(147)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(147)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(147) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(147) is a control-delay.
    cp_element_147_delay: control_delay_element  generic map(name => " 147_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(145), ack => access_T_CP_0_elements(147), clk => clk, reset =>reset);
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	152 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	153 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/addr_of_133_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/addr_of_133_request/$entry
      -- CP-element group 148: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/addr_of_133_request/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(148)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(148)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(148) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:addr_of_133_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(148), ack => addr_of_133_final_reg_req_0); -- 
    access_T_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(152) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	9 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	157 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	154 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/addr_of_133_update_start_
      -- CP-element group 149: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/addr_of_133_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/addr_of_133_complete/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(149)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(149)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(149) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:addr_of_133_final_reg_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(149), ack => addr_of_133_final_reg_req_1); -- 
    access_T_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	9 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	153 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_final_index_sum_regn_update_start
      -- CP-element group 150: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_final_index_sum_regn_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_final_index_sum_regn_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(150)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(150)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(150) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:array_obj_ref_132_index_offset_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(150), ack => array_obj_ref_132_index_offset_req_1); -- 
    access_T_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	18 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	204 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	16 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_final_index_sum_regn_sample_complete
      -- CP-element group 151: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_final_index_sum_regn_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(151)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(151)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(151) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:array_obj_ref_132_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_132_index_offset_ack_0, ack => access_T_CP_0_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	148 
    -- CP-element group 152:  members (8) 
      -- CP-element group 152: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_root_address_calculated
      -- CP-element group 152: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_offset_calculated
      -- CP-element group 152: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_final_index_sum_regn_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_final_index_sum_regn_Update/ack
      -- CP-element group 152: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_base_plus_offset/$entry
      -- CP-element group 152: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_base_plus_offset/$exit
      -- CP-element group 152: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_base_plus_offset/sum_rename_req
      -- CP-element group 152: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/array_obj_ref_132_base_plus_offset/sum_rename_ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(152)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(152)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(152) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:array_obj_ref_132_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_132_index_offset_ack_1, ack => access_T_CP_0_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: 	150 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/addr_of_133_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/addr_of_133_request/$exit
      -- CP-element group 153: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/addr_of_133_request/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(153)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(153)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(153) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:addr_of_133_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_133_final_reg_ack_0, ack => access_T_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	149 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (19) 
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/addr_of_133_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/addr_of_133_complete/$exit
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/addr_of_133_complete/ack
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(154)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(154)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(154) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:addr_of_133_final_reg_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_133_final_reg_ack_1, ack => access_T_CP_0_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (5) 
      -- CP-element group 155: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Sample/word_access_start/$entry
      -- CP-element group 155: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Sample/word_access_start/word_0/$entry
      -- CP-element group 155: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group access_T_CP_0_elements(155)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(155)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(155) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:ptr_deref_137_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(155), ack => ptr_deref_137_load_0_req_0); -- 
    access_T_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(154) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	165 
    -- CP-element group 156: 	169 
    -- CP-element group 156: 	173 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_update_start_
      -- CP-element group 156: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Update/word_access_complete/$entry
      -- CP-element group 156: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Update/word_access_complete/word_0/$entry
      -- CP-element group 156: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group access_T_CP_0_elements(156)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(156)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(156) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:ptr_deref_137_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(156), ack => ptr_deref_137_load_0_req_1); -- 
    access_T_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(161) & access_T_CP_0_elements(165) & access_T_CP_0_elements(169) & access_T_CP_0_elements(173);
      gj_access_T_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	149 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (5) 
      -- CP-element group 157: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Sample/word_access_start/$exit
      -- CP-element group 157: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Sample/word_access_start/word_0/$exit
      -- CP-element group 157: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group access_T_CP_0_elements(157)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(157)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(157) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:ptr_deref_137_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_137_load_0_ack_0, ack => access_T_CP_0_elements(157)); -- 
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	163 
    -- CP-element group 158: 	167 
    -- CP-element group 158: 	171 
    -- CP-element group 158:  members (9) 
      -- CP-element group 158: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Update/word_access_complete/$exit
      -- CP-element group 158: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Update/word_access_complete/word_0/$exit
      -- CP-element group 158: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Update/word_access_complete/word_0/ca
      -- CP-element group 158: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Update/ptr_deref_137_Merge/$entry
      -- CP-element group 158: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Update/ptr_deref_137_Merge/$exit
      -- CP-element group 158: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Update/ptr_deref_137_Merge/merge_req
      -- CP-element group 158: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/ptr_deref_137_Update/ptr_deref_137_Merge/merge_ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(158)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(158)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(158) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:ptr_deref_137_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_137_load_0_ack_1, ack => access_T_CP_0_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_141_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_141_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_141_Sample/rr
      -- 
    -- logger for CP element group access_T_CP_0_elements(159)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(159)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(159) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_141_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(159), ack => slice_141_inst_req_0); -- 
    access_T_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(161);
      gj_access_T_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	180 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_141_update_start_
      -- CP-element group 160: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_141_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_141_Update/cr
      -- 
    -- logger for CP element group access_T_CP_0_elements(160)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(160)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(160) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_141_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(160), ack => slice_141_inst_req_1); -- 
    access_T_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	159 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_141_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_141_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_141_Sample/ra
      -- 
    -- logger for CP element group access_T_CP_0_elements(161)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(161)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(161) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_141_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_141_inst_ack_0, ack => access_T_CP_0_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	179 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_141_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_141_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_141_Update/ca
      -- 
    -- logger for CP element group access_T_CP_0_elements(162)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(162)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(162) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_141_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_141_inst_ack_1, ack => access_T_CP_0_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	158 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_145_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_145_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_145_Sample/rr
      -- 
    -- logger for CP element group access_T_CP_0_elements(163)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(163)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(163) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_145_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(163), ack => slice_145_inst_req_0); -- 
    access_T_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(165);
      gj_access_T_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	187 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_145_update_start_
      -- CP-element group 164: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_145_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_145_Update/cr
      -- 
    -- logger for CP element group access_T_CP_0_elements(164)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(164)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(164) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_145_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(164), ack => slice_145_inst_req_1); -- 
    access_T_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	156 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_145_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_145_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_145_Sample/ra
      -- 
    -- logger for CP element group access_T_CP_0_elements(165)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(165)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(165) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_145_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_145_inst_ack_0, ack => access_T_CP_0_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	186 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_145_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_145_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_145_Update/ca
      -- 
    -- logger for CP element group access_T_CP_0_elements(166)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(166)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(166) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_145_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_145_inst_ack_1, ack => access_T_CP_0_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	158 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_149_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_149_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_149_Sample/rr
      -- 
    -- logger for CP element group access_T_CP_0_elements(167)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(167)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(167) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_149_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(167), ack => slice_149_inst_req_0); -- 
    access_T_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(169);
      gj_access_T_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	194 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_149_update_start_
      -- CP-element group 168: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_149_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_149_Update/cr
      -- 
    -- logger for CP element group access_T_CP_0_elements(168)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(168)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(168) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_149_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(168), ack => slice_149_inst_req_1); -- 
    access_T_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	156 
    -- CP-element group 169: 	167 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_149_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_149_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_149_Sample/ra
      -- 
    -- logger for CP element group access_T_CP_0_elements(169)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(169)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(169) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_149_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_149_inst_ack_0, ack => access_T_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	193 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_149_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_149_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_149_Update/ca
      -- 
    -- logger for CP element group access_T_CP_0_elements(170)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(170)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(170) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_149_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_149_inst_ack_1, ack => access_T_CP_0_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	158 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_153_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_153_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_153_Sample/rr
      -- 
    -- logger for CP element group access_T_CP_0_elements(171)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(171)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(171) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_153_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(171), ack => slice_153_inst_req_0); -- 
    access_T_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(173);
      gj_access_T_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	201 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_153_update_start_
      -- CP-element group 172: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_153_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_153_Update/cr
      -- 
    -- logger for CP element group access_T_CP_0_elements(172)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(172)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(172) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_153_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(172), ack => slice_153_inst_req_1); -- 
    access_T_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	156 
    -- CP-element group 173: 	171 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_153_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_153_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_153_Sample/ra
      -- 
    -- logger for CP element group access_T_CP_0_elements(173)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(173)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(173) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_153_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_153_inst_ack_0, ack => access_T_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	200 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_153_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_153_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/slice_153_Update/ca
      -- 
    -- logger for CP element group access_T_CP_0_elements(174)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(174)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(174) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:slice_153_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_153_inst_ack_1, ack => access_T_CP_0_elements(174)); -- 
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	37 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_157_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_157_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_157_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(175)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(175)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(175) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c1_155_delayed_14_0_155_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(175), ack => W_c1_155_delayed_14_0_155_inst_req_0); -- 
    access_T_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(37) & access_T_CP_0_elements(177);
      gj_access_T_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	180 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_157_update_start_
      -- CP-element group 176: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_157_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_157_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(176)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(176)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(176) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c1_155_delayed_14_0_155_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(176), ack => W_c1_155_delayed_14_0_155_inst_req_1); -- 
    access_T_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	33 
    -- CP-element group 177: 	175 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_157_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_157_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_157_Sample/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(177)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(177)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(177) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c1_155_delayed_14_0_155_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_155_delayed_14_0_155_inst_ack_0, ack => access_T_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_157_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_157_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_157_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(178)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(178)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(178) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c1_155_delayed_14_0_155_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_155_delayed_14_0_155_inst_ack_1, ack => access_T_CP_0_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	162 
    -- CP-element group 179: 	178 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	202 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_159_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_159_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_159_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(179)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(179)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(179) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_159_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(179), ack => WPIPE_input_pipe1_159_inst_req_0); -- 
    access_T_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(162) & access_T_CP_0_elements(178) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	160 
    -- CP-element group 180: 	176 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_159_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_159_update_start_
      -- CP-element group 180: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_159_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_159_Sample/ack
      -- CP-element group 180: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_159_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_159_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(180)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(180)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(180) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_159_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_159_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_159_inst_ack_0, ack => access_T_CP_0_elements(180)); -- 
    req_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(180), ack => WPIPE_input_pipe1_159_inst_req_1); -- 
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	186 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_159_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_159_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_159_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(181)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(181)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(181) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_159_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_159_inst_ack_1, ack => access_T_CP_0_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	37 
    -- CP-element group 182: 	75 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_164_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_164_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_164_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(182)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(182)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(182) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c2_159_delayed_14_0_162_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(182), ack => W_c2_159_delayed_14_0_162_inst_req_0); -- 
    access_T_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(37) & access_T_CP_0_elements(75) & access_T_CP_0_elements(184);
      gj_access_T_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	187 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_164_update_start_
      -- CP-element group 183: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_164_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_164_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(183)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(183)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(183) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c2_159_delayed_14_0_162_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(183), ack => W_c2_159_delayed_14_0_162_inst_req_1); -- 
    access_T_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	33 
    -- CP-element group 184: 	71 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_164_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_164_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_164_Sample/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(184)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(184)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(184) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c2_159_delayed_14_0_162_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_159_delayed_14_0_162_inst_ack_0, ack => access_T_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_164_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_164_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_164_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(185)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(185)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(185) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c2_159_delayed_14_0_162_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_159_delayed_14_0_162_inst_ack_1, ack => access_T_CP_0_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	166 
    -- CP-element group 186: 	181 
    -- CP-element group 186: 	185 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_166_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_166_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_166_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(186)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(186)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(186) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_166_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(186), ack => WPIPE_input_pipe1_166_inst_req_0); -- 
    access_T_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(166) & access_T_CP_0_elements(181) & access_T_CP_0_elements(185) & access_T_CP_0_elements(188);
      gj_access_T_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	164 
    -- CP-element group 187: 	183 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_166_Sample/ack
      -- CP-element group 187: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_166_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_166_Update/req
      -- CP-element group 187: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_166_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_166_update_start_
      -- CP-element group 187: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_166_Sample/$exit
      -- 
    -- logger for CP element group access_T_CP_0_elements(187)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(187)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(187) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_166_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_166_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_166_inst_ack_0, ack => access_T_CP_0_elements(187)); -- 
    req_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(187), ack => WPIPE_input_pipe1_166_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	193 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_166_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_166_Update/ack
      -- CP-element group 188: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_166_update_completed_
      -- 
    -- logger for CP element group access_T_CP_0_elements(188)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(188)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(188) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_166_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_166_inst_ack_1, ack => access_T_CP_0_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	37 
    -- CP-element group 189: 	75 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_171_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_171_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_171_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(189)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(189)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(189) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c3_163_delayed_14_0_169_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(189), ack => W_c3_163_delayed_14_0_169_inst_req_0); -- 
    access_T_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(37) & access_T_CP_0_elements(75) & access_T_CP_0_elements(191);
      gj_access_T_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	194 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_171_update_start_
      -- CP-element group 190: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_171_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_171_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(190)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(190)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(190) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c3_163_delayed_14_0_169_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(190), ack => W_c3_163_delayed_14_0_169_inst_req_1); -- 
    access_T_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	33 
    -- CP-element group 191: 	71 
    -- CP-element group 191: 	189 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_171_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_171_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_171_Sample/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(191)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(191)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(191) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c3_163_delayed_14_0_169_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_163_delayed_14_0_169_inst_ack_0, ack => access_T_CP_0_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_171_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_171_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_171_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(192)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(192)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(192) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c3_163_delayed_14_0_169_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_163_delayed_14_0_169_inst_ack_1, ack => access_T_CP_0_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	170 
    -- CP-element group 193: 	188 
    -- CP-element group 193: 	192 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_173_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_173_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_173_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(193)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(193)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(193) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_173_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(193), ack => WPIPE_input_pipe1_173_inst_req_0); -- 
    access_T_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(170) & access_T_CP_0_elements(188) & access_T_CP_0_elements(192) & access_T_CP_0_elements(195);
      gj_access_T_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	168 
    -- CP-element group 194: 	190 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_173_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_173_update_start_
      -- CP-element group 194: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_173_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_173_Sample/ack
      -- CP-element group 194: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_173_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_173_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(194)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(194)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(194) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_173_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_173_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_173_inst_ack_0, ack => access_T_CP_0_elements(194)); -- 
    req_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(194), ack => WPIPE_input_pipe1_173_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	200 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_173_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_173_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_173_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(195)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(195)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(195) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_173_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_173_inst_ack_1, ack => access_T_CP_0_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	37 
    -- CP-element group 196: 	75 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_178_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_178_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_178_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(196)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(196)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(196) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c4_167_delayed_14_0_176_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(196), ack => W_c4_167_delayed_14_0_176_inst_req_0); -- 
    access_T_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(37) & access_T_CP_0_elements(75) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	201 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_178_update_start_
      -- CP-element group 197: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_178_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_178_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(197)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(197)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(197) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c4_167_delayed_14_0_176_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(197), ack => W_c4_167_delayed_14_0_176_inst_req_1); -- 
    access_T_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	33 
    -- CP-element group 198: 	71 
    -- CP-element group 198: 	196 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_178_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_178_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_178_Sample/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(198)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(198)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(198) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c4_167_delayed_14_0_176_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_167_delayed_14_0_176_inst_ack_0, ack => access_T_CP_0_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_178_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_178_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/assign_stmt_178_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(199)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(199)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(199) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:W_c4_167_delayed_14_0_176_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_167_delayed_14_0_176_inst_ack_1, ack => access_T_CP_0_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	174 
    -- CP-element group 200: 	195 
    -- CP-element group 200: 	199 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_180_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_180_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_180_Sample/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(200)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(200)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(200) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_180_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(200), ack => WPIPE_input_pipe1_180_inst_req_0); -- 
    access_T_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(174) & access_T_CP_0_elements(195) & access_T_CP_0_elements(199) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	172 
    -- CP-element group 201: 	197 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_180_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_180_update_start_
      -- CP-element group 201: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_180_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_180_Sample/ack
      -- CP-element group 201: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_180_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_180_Update/req
      -- 
    -- logger for CP element group access_T_CP_0_elements(201)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(201)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(201) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_180_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_180_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_180_inst_ack_0, ack => access_T_CP_0_elements(201)); -- 
    req_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(201), ack => WPIPE_input_pipe1_180_inst_req_1); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	179 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_180_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_180_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/WPIPE_input_pipe1_180_Update/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(202)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(202)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(202) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:WPIPE_input_pipe1_180_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_180_inst_ack_1, ack => access_T_CP_0_elements(202)); -- 
    -- CP-element group 203:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	9 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	10 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group access_T_CP_0_elements(203)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(203)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(203) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group access_T_CP_0_elements(203) is a control-delay.
    cp_element_203_delay: control_delay_element  generic map(name => " 203_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(9), ack => access_T_CP_0_elements(203), clk => clk, reset =>reset);
    -- CP-element group 204:  join  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	12 
    -- CP-element group 204: 	151 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	6 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_25/do_while_stmt_43/do_while_stmt_43_loop_body/$exit
      -- 
    -- logger for CP element group access_T_CP_0_elements(204)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(204)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(204) fired."); 
        -- 
      end if; --
    end process; 
    access_T_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(12) & access_T_CP_0_elements(151) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	5 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_25/do_while_stmt_43/loop_exit/$exit
      -- CP-element group 205: 	 branch_block_stmt_25/do_while_stmt_43/loop_exit/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(205)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(205)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(205) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:do_while_stmt_43_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_43_branch_ack_0, ack => access_T_CP_0_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	5 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (2) 
      -- CP-element group 206: 	 branch_block_stmt_25/do_while_stmt_43/loop_taken/$exit
      -- CP-element group 206: 	 branch_block_stmt_25/do_while_stmt_43/loop_taken/ack
      -- 
    -- logger for CP element group access_T_CP_0_elements(206)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(206)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(206) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:do_while_stmt_43_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_43_branch_ack_1, ack => access_T_CP_0_elements(206)); -- 
    -- CP-element group 207:  transition  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	3 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	1 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_25/do_while_stmt_43/$exit
      -- 
    -- logger for CP element group access_T_CP_0_elements(207)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and access_T_CP_0_elements(207)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:access_T:CP:access_T_CP_0_elements(207) fired."); 
        -- 
      end if; --
    end process; 
    access_T_CP_0_elements(207) <= access_T_CP_0_elements(3);
    access_T_do_while_stmt_43_terminator_636: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_43_terminator_636", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(6),loop_continue => access_T_CP_0_elements(206),loop_terminate => access_T_CP_0_elements(205),loop_back => access_T_CP_0_elements(4),loop_exit => access_T_CP_0_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_45_phi_seq_78_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(19);
      access_T_CP_0_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(26);
      access_T_CP_0_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(27);
      access_T_CP_0_elements(20) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(21);
      access_T_CP_0_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(28);
      access_T_CP_0_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(30);
      access_T_CP_0_elements(22) <= phi_mux_reqs(1);
      phi_stmt_45_phi_seq_78 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_45_phi_seq_78") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(11), 
          phi_sample_ack => access_T_CP_0_elements(17), 
          phi_update_req => access_T_CP_0_elements(13), 
          phi_update_ack => access_T_CP_0_elements(18), 
          phi_mux_ack => access_T_CP_0_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_50_phi_seq_122_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(38);
      access_T_CP_0_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(45);
      access_T_CP_0_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(46);
      access_T_CP_0_elements(39) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(40);
      access_T_CP_0_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(47);
      access_T_CP_0_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(49);
      access_T_CP_0_elements(41) <= phi_mux_reqs(1);
      phi_stmt_50_phi_seq_122 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_50_phi_seq_122") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(34), 
          phi_sample_ack => access_T_CP_0_elements(35), 
          phi_update_req => access_T_CP_0_elements(36), 
          phi_update_ack => access_T_CP_0_elements(37), 
          phi_mux_ack => access_T_CP_0_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_56_phi_seq_176_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(59);
      access_T_CP_0_elements(62)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(64);
      access_T_CP_0_elements(63)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(65);
      access_T_CP_0_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(57);
      access_T_CP_0_elements(66)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(68);
      access_T_CP_0_elements(67)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(69);
      access_T_CP_0_elements(58) <= phi_mux_reqs(1);
      phi_stmt_56_phi_seq_176 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_56_phi_seq_176") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(53), 
          phi_sample_ack => access_T_CP_0_elements(54), 
          phi_update_req => access_T_CP_0_elements(55), 
          phi_update_ack => access_T_CP_0_elements(56), 
          phi_mux_ack => access_T_CP_0_elements(61), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_60_phi_seq_230_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(76);
      access_T_CP_0_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(83);
      access_T_CP_0_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(84);
      access_T_CP_0_elements(77) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(78);
      access_T_CP_0_elements(85)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(89);
      access_T_CP_0_elements(86)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(90);
      access_T_CP_0_elements(79) <= phi_mux_reqs(1);
      phi_stmt_60_phi_seq_230 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_60_phi_seq_230") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(72), 
          phi_sample_ack => access_T_CP_0_elements(73), 
          phi_update_req => access_T_CP_0_elements(74), 
          phi_update_ack => access_T_CP_0_elements(75), 
          phi_mux_ack => access_T_CP_0_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_65_phi_seq_274_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(99);
      access_T_CP_0_elements(102)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(102);
      access_T_CP_0_elements(103)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(104);
      access_T_CP_0_elements(100) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(97);
      access_T_CP_0_elements(106)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(108);
      access_T_CP_0_elements(107)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(109);
      access_T_CP_0_elements(98) <= phi_mux_reqs(1);
      phi_stmt_65_phi_seq_274 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_65_phi_seq_274") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(93), 
          phi_sample_ack => access_T_CP_0_elements(94), 
          phi_update_req => access_T_CP_0_elements(95), 
          phi_update_ack => access_T_CP_0_elements(96), 
          phi_mux_ack => access_T_CP_0_elements(101), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_70_phi_seq_318_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(118);
      access_T_CP_0_elements(121)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(121);
      access_T_CP_0_elements(122)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(123);
      access_T_CP_0_elements(119) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(116);
      access_T_CP_0_elements(125)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(127);
      access_T_CP_0_elements(126)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(128);
      access_T_CP_0_elements(117) <= phi_mux_reqs(1);
      phi_stmt_70_phi_seq_318 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_70_phi_seq_318") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(112), 
          phi_sample_ack => access_T_CP_0_elements(113), 
          phi_update_req => access_T_CP_0_elements(114), 
          phi_update_ack => access_T_CP_0_elements(115), 
          phi_mux_ack => access_T_CP_0_elements(120), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_75_phi_seq_362_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(135);
      access_T_CP_0_elements(140)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(142);
      access_T_CP_0_elements(141)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(143);
      access_T_CP_0_elements(136) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(137);
      access_T_CP_0_elements(144)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(144);
      access_T_CP_0_elements(145)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(146);
      access_T_CP_0_elements(138) <= phi_mux_reqs(1);
      phi_stmt_75_phi_seq_362 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_75_phi_seq_362") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(131), 
          phi_sample_ack => access_T_CP_0_elements(132), 
          phi_update_req => access_T_CP_0_elements(133), 
          phi_update_ack => access_T_CP_0_elements(134), 
          phi_mux_ack => access_T_CP_0_elements(139), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_30_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(7);
        preds(1)  <= access_T_CP_0_elements(8);
        entry_tmerge_30 : transition_merge -- 
          generic map(name => " entry_tmerge_30")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_124_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_204_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_217_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_230_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_240_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_292_wire : std_logic_vector(15 downto 0);
    signal ADD_u64_u64_277_wire : std_logic_vector(63 downto 0);
    signal AND_u1_u1_106_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_113_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_212_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_226_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_227_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_93_wire : std_logic_vector(0 downto 0);
    signal AND_u32_u32_259_wire : std_logic_vector(31 downto 0);
    signal EQ_u2_u1_102_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_109_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_116_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_89_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_96_wire : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_273_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_239_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_241_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_29_wire : std_logic_vector(15 downto 0);
    signal MUL_u32_u32_248_wire : std_logic_vector(31 downto 0);
    signal MUX_205_wire : std_logic_vector(15 downto 0);
    signal MUX_218_wire : std_logic_vector(15 downto 0);
    signal MUX_299_wire : std_logic_vector(15 downto 0);
    signal MUX_305_wire : std_logic_vector(15 downto 0);
    signal NEQ_u16_u1_311_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_117_wire : std_logic_vector(0 downto 0);
    signal R_address_131_resized : std_logic_vector(13 downto 0);
    signal R_address_131_scaled : std_logic_vector(13 downto 0);
    signal SUB_u16_u16_285_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_297_wire : std_logic_vector(15 downto 0);
    signal UGT_u16_u1_105_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_112_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_294_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_92_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_302_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_38_wire : std_logic_vector(0 downto 0);
    signal address_45 : std_logic_vector(63 downto 0);
    signal array_obj_ref_132_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_132_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_132_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_132_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_132_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_132_root_address : std_logic_vector(13 downto 0);
    signal c1_155_delayed_14_0_157 : std_logic_vector(0 downto 0);
    signal c1_85 : std_logic_vector(0 downto 0);
    signal c2_159_delayed_14_0_164 : std_logic_vector(0 downto 0);
    signal c2_98 : std_logic_vector(0 downto 0);
    signal c3_119 : std_logic_vector(0 downto 0);
    signal c3_163_delayed_14_0_171 : std_logic_vector(0 downto 0);
    signal c4_127 : std_logic_vector(0 downto 0);
    signal c4_167_delayed_14_0_178 : std_logic_vector(0 downto 0);
    signal col_70 : std_logic_vector(15 downto 0);
    signal col_done_197 : std_logic_vector(0 downto 0);
    signal fetch_addr_134 : std_logic_vector(31 downto 0);
    signal flag1_187 : std_logic_vector(0 downto 0);
    signal fn_blk_42 : std_logic_vector(15 downto 0);
    signal konst_101_wire_constant : std_logic_vector(1 downto 0);
    signal konst_104_wire_constant : std_logic_vector(15 downto 0);
    signal konst_108_wire_constant : std_logic_vector(1 downto 0);
    signal konst_111_wire_constant : std_logic_vector(15 downto 0);
    signal konst_115_wire_constant : std_logic_vector(1 downto 0);
    signal konst_125_wire_constant : std_logic_vector(15 downto 0);
    signal konst_201_wire_constant : std_logic_vector(15 downto 0);
    signal konst_203_wire_constant : std_logic_vector(15 downto 0);
    signal konst_214_wire_constant : std_logic_vector(15 downto 0);
    signal konst_216_wire_constant : std_logic_vector(15 downto 0);
    signal konst_229_wire_constant : std_logic_vector(15 downto 0);
    signal konst_258_wire_constant : std_logic_vector(31 downto 0);
    signal konst_266_wire_constant : std_logic_vector(1 downto 0);
    signal konst_272_wire_constant : std_logic_vector(31 downto 0);
    signal konst_276_wire_constant : std_logic_vector(63 downto 0);
    signal konst_293_wire_constant : std_logic_vector(15 downto 0);
    signal konst_295_wire_constant : std_logic_vector(15 downto 0);
    signal konst_301_wire_constant : std_logic_vector(15 downto 0);
    signal konst_304_wire_constant : std_logic_vector(15 downto 0);
    signal konst_37_wire_constant : std_logic_vector(15 downto 0);
    signal konst_40_wire_constant : std_logic_vector(15 downto 0);
    signal konst_83_wire_constant : std_logic_vector(1 downto 0);
    signal konst_88_wire_constant : std_logic_vector(1 downto 0);
    signal konst_91_wire_constant : std_logic_vector(15 downto 0);
    signal konst_95_wire_constant : std_logic_vector(1 downto 0);
    signal m_factor_31 : std_logic_vector(31 downto 0);
    signal n_address_279 : std_logic_vector(63 downto 0);
    signal n_address_279_47_buffered : std_logic_vector(63 downto 0);
    signal n_blk_307 : std_logic_vector(15 downto 0);
    signal n_blk_307_62_buffered : std_logic_vector(15 downto 0);
    signal n_col_221 : std_logic_vector(15 downto 0);
    signal n_col_221_74_buffered : std_logic_vector(15 downto 0);
    signal n_left_287 : std_logic_vector(15 downto 0);
    signal n_left_287_59_buffered : std_logic_vector(15 downto 0);
    signal n_row_233 : std_logic_vector(15 downto 0);
    signal n_row_233_77_buffered : std_logic_vector(15 downto 0);
    signal n_winr_208 : std_logic_vector(15 downto 0);
    signal n_winr_208_69_buffered : std_logic_vector(15 downto 0);
    signal n_word_start_268 : std_logic_vector(1 downto 0);
    signal n_word_start_268_52_buffered : std_logic_vector(1 downto 0);
    signal na1_243 : std_logic_vector(31 downto 0);
    signal na2_250 : std_logic_vector(31 downto 0);
    signal na3_255 : std_logic_vector(31 downto 0);
    signal na4_261 : std_logic_vector(15 downto 0);
    signal nl_start_34 : std_logic_vector(15 downto 0);
    signal nl_start_34_58_buffered : std_logic_vector(15 downto 0);
    signal num_blk_60 : std_logic_vector(15 downto 0);
    signal num_left_56 : std_logic_vector(15 downto 0);
    signal ptr_deref_137_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_137_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_137_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_137_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_137_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_75 : std_logic_vector(15 downto 0);
    signal type_cast_123_wire : std_logic_vector(15 downto 0);
    signal type_cast_247_wire : std_logic_vector(31 downto 0);
    signal type_cast_265_wire : std_logic_vector(1 downto 0);
    signal type_cast_274_wire : std_logic_vector(63 downto 0);
    signal type_cast_49_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_55_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_64_wire : std_logic_vector(15 downto 0);
    signal type_cast_68_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_73_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_79_wire_constant : std_logic_vector(15 downto 0);
    signal w1_142 : std_logic_vector(15 downto 0);
    signal w2_146 : std_logic_vector(15 downto 0);
    signal w3_150 : std_logic_vector(15 downto 0);
    signal w4_154 : std_logic_vector(15 downto 0);
    signal winr_65 : std_logic_vector(15 downto 0);
    signal winr_done_192 : std_logic_vector(0 downto 0);
    signal word_read_138 : std_logic_vector(63 downto 0);
    signal word_start_50 : std_logic_vector(1 downto 0);
    -- 
  begin -- 
    array_obj_ref_132_constant_part_of_offset <= "00000000000000";
    array_obj_ref_132_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_132_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_132_resized_base_address <= "00000000000000";
    konst_101_wire_constant <= "00";
    konst_104_wire_constant <= "0000000000000010";
    konst_108_wire_constant <= "01";
    konst_111_wire_constant <= "0000000000000001";
    konst_115_wire_constant <= "10";
    konst_125_wire_constant <= "0000000000000011";
    konst_201_wire_constant <= "0000000000000000";
    konst_203_wire_constant <= "0000000000000001";
    konst_214_wire_constant <= "0000000000000000";
    konst_216_wire_constant <= "0000000000000001";
    konst_229_wire_constant <= "0000000000000001";
    konst_258_wire_constant <= "00000000000000000000000000000011";
    konst_266_wire_constant <= "00";
    konst_272_wire_constant <= "00000000000000000000000000000010";
    konst_276_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_293_wire_constant <= "0000000000000100";
    konst_295_wire_constant <= "0000000000000100";
    konst_301_wire_constant <= "0000000000000100";
    konst_304_wire_constant <= "0000000000000100";
    konst_37_wire_constant <= "0000000000000100";
    konst_40_wire_constant <= "0000000000000100";
    konst_83_wire_constant <= "00";
    konst_88_wire_constant <= "00";
    konst_91_wire_constant <= "0000000000000001";
    konst_95_wire_constant <= "01";
    ptr_deref_137_word_offset_0 <= "00000000000000";
    type_cast_49_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_55_wire_constant <= "00";
    type_cast_68_wire_constant <= "0000000000000000";
    type_cast_73_wire_constant <= "0000000000000000";
    type_cast_79_wire_constant <= "0000000000000000";
    -- logger for phi phi_stmt_45
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_45_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_45:input-0 n_address_279_47_buffered= " & Convert_SLV_To_Hex_String(n_address_279_47_buffered));
          --
        end if;
        if phi_stmt_45_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_45:input-1 type_cast_49_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_49_wire_constant));
          --
        end if;
        if phi_stmt_45_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:access_T:DP:phi_stmt_45:sample-completed");
          --
        end if;
        if phi_stmt_45_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:access_T:DP:phi_stmt_45:output address_45= " & Convert_SLV_To_Hex_String(address_45));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_45: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_address_279_47_buffered & type_cast_49_wire_constant;
      req <= phi_stmt_45_req_0 & phi_stmt_45_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_45",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_45_ack_0,
          idata => idata,
          odata => address_45,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_45
    -- logger for phi phi_stmt_50
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_50_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_50:input-0 n_word_start_268_52_buffered= " & Convert_SLV_To_Hex_String(n_word_start_268_52_buffered));
          --
        end if;
        if phi_stmt_50_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_50:input-1 type_cast_55_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_55_wire_constant));
          --
        end if;
        if phi_stmt_50_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:access_T:DP:phi_stmt_50:sample-completed");
          --
        end if;
        if phi_stmt_50_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:access_T:DP:phi_stmt_50:output word_start_50= " & Convert_SLV_To_Hex_String(word_start_50));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_50: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_word_start_268_52_buffered & type_cast_55_wire_constant;
      req <= phi_stmt_50_req_0 & phi_stmt_50_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_50",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_50_ack_0,
          idata => idata,
          odata => word_start_50,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_50
    -- logger for phi phi_stmt_56
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_56_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_56:input-0 nl_start_34_58_buffered= " & Convert_SLV_To_Hex_String(nl_start_34_58_buffered));
          --
        end if;
        if phi_stmt_56_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_56:input-1 n_left_287_59_buffered= " & Convert_SLV_To_Hex_String(n_left_287_59_buffered));
          --
        end if;
        if phi_stmt_56_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:access_T:DP:phi_stmt_56:sample-completed");
          --
        end if;
        if phi_stmt_56_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:access_T:DP:phi_stmt_56:output num_left_56= " & Convert_SLV_To_Hex_String(num_left_56));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_56: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nl_start_34_58_buffered & n_left_287_59_buffered;
      req <= phi_stmt_56_req_0 & phi_stmt_56_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_56",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_56_ack_0,
          idata => idata,
          odata => num_left_56,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_56
    -- logger for phi phi_stmt_60
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_60_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_60:input-0 n_blk_307_62_buffered= " & Convert_SLV_To_Hex_String(n_blk_307_62_buffered));
          --
        end if;
        if phi_stmt_60_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_60:input-1 type_cast_64_wire= " & Convert_SLV_To_Hex_String(type_cast_64_wire));
          --
        end if;
        if phi_stmt_60_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:access_T:DP:phi_stmt_60:sample-completed");
          --
        end if;
        if phi_stmt_60_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:access_T:DP:phi_stmt_60:output num_blk_60= " & Convert_SLV_To_Hex_String(num_blk_60));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_60: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_blk_307_62_buffered & type_cast_64_wire;
      req <= phi_stmt_60_req_0 & phi_stmt_60_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_60",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_60_ack_0,
          idata => idata,
          odata => num_blk_60,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_60
    -- logger for phi phi_stmt_65
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_65_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_65:input-0 type_cast_68_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_68_wire_constant));
          --
        end if;
        if phi_stmt_65_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_65:input-1 n_winr_208_69_buffered= " & Convert_SLV_To_Hex_String(n_winr_208_69_buffered));
          --
        end if;
        if phi_stmt_65_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:access_T:DP:phi_stmt_65:sample-completed");
          --
        end if;
        if phi_stmt_65_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:access_T:DP:phi_stmt_65:output winr_65= " & Convert_SLV_To_Hex_String(winr_65));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_65: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_68_wire_constant & n_winr_208_69_buffered;
      req <= phi_stmt_65_req_0 & phi_stmt_65_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_65",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_65_ack_0,
          idata => idata,
          odata => winr_65,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_65
    -- logger for phi phi_stmt_70
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_70_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_70:input-0 type_cast_73_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_73_wire_constant));
          --
        end if;
        if phi_stmt_70_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_70:input-1 n_col_221_74_buffered= " & Convert_SLV_To_Hex_String(n_col_221_74_buffered));
          --
        end if;
        if phi_stmt_70_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:access_T:DP:phi_stmt_70:sample-completed");
          --
        end if;
        if phi_stmt_70_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:access_T:DP:phi_stmt_70:output col_70= " & Convert_SLV_To_Hex_String(col_70));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_70: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_73_wire_constant & n_col_221_74_buffered;
      req <= phi_stmt_70_req_0 & phi_stmt_70_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_70",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_70_ack_0,
          idata => idata,
          odata => col_70,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_70
    -- logger for phi phi_stmt_75
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_75_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_75:input-0 n_row_233_77_buffered= " & Convert_SLV_To_Hex_String(n_row_233_77_buffered));
          --
        end if;
        if phi_stmt_75_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:access_T:DP:phi_stmt_75:input-1 type_cast_79_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_79_wire_constant));
          --
        end if;
        if phi_stmt_75_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:access_T:DP:phi_stmt_75:sample-completed");
          --
        end if;
        if phi_stmt_75_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:access_T:DP:phi_stmt_75:output row_75= " & Convert_SLV_To_Hex_String(row_75));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_75: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_row_233_77_buffered & type_cast_79_wire_constant;
      req <= phi_stmt_75_req_0 & phi_stmt_75_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_75",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_75_ack_0,
          idata => idata,
          odata => row_75,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_75
    -- logger for split-operator MUX_205_inst flow-through 
    process(MUX_205_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUX_205_inst:flowthrough inputs: " & " winr_done_192 = "& Convert_SLV_To_Hex_String(winr_done_192) & " konst_201_wire_constant = "& Convert_SLV_To_Hex_String(konst_201_wire_constant) & " ADD_u16_u16_204_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_204_wire) & " outputs:" & " MUX_205_wire= "  & Convert_SLV_To_Hex_String(MUX_205_wire));
      --
    end process; 
    -- flow-through select operator MUX_205_inst
    MUX_205_wire <= konst_201_wire_constant when (winr_done_192(0) /=  '0') else ADD_u16_u16_204_wire;
    -- logger for split-operator MUX_207_inst flow-through 
    process(n_winr_208) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUX_207_inst:flowthrough inputs: " & " flag1_187 = "& Convert_SLV_To_Hex_String(flag1_187) & " MUX_205_wire = "& Convert_SLV_To_Hex_String(MUX_205_wire) & " winr_65 = "& Convert_SLV_To_Hex_String(winr_65) & " outputs:" & " n_winr_208= "  & Convert_SLV_To_Hex_String(n_winr_208));
      --
    end process; 
    -- flow-through select operator MUX_207_inst
    n_winr_208 <= MUX_205_wire when (flag1_187(0) /=  '0') else winr_65;
    -- logger for split-operator MUX_218_inst flow-through 
    process(MUX_218_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUX_218_inst:flowthrough inputs: " & " col_done_197 = "& Convert_SLV_To_Hex_String(col_done_197) & " konst_214_wire_constant = "& Convert_SLV_To_Hex_String(konst_214_wire_constant) & " ADD_u16_u16_217_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_217_wire) & " outputs:" & " MUX_218_wire= "  & Convert_SLV_To_Hex_String(MUX_218_wire));
      --
    end process; 
    -- flow-through select operator MUX_218_inst
    MUX_218_wire <= konst_214_wire_constant when (col_done_197(0) /=  '0') else ADD_u16_u16_217_wire;
    -- logger for split-operator MUX_220_inst flow-through 
    process(n_col_221) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUX_220_inst:flowthrough inputs: " & " AND_u1_u1_212_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_212_wire) & " MUX_218_wire = "& Convert_SLV_To_Hex_String(MUX_218_wire) & " col_70 = "& Convert_SLV_To_Hex_String(col_70) & " outputs:" & " n_col_221= "  & Convert_SLV_To_Hex_String(n_col_221));
      --
    end process; 
    -- flow-through select operator MUX_220_inst
    n_col_221 <= MUX_218_wire when (AND_u1_u1_212_wire(0) /=  '0') else col_70;
    -- logger for split-operator MUX_232_inst flow-through 
    process(n_row_233) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUX_232_inst:flowthrough inputs: " & " AND_u1_u1_227_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_227_wire) & " ADD_u16_u16_230_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_230_wire) & " row_75 = "& Convert_SLV_To_Hex_String(row_75) & " outputs:" & " n_row_233= "  & Convert_SLV_To_Hex_String(n_row_233));
      --
    end process; 
    -- flow-through select operator MUX_232_inst
    n_row_233 <= ADD_u16_u16_230_wire when (AND_u1_u1_227_wire(0) /=  '0') else row_75;
    -- logger for split-operator MUX_267_inst flow-through 
    process(n_word_start_268) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUX_267_inst:flowthrough inputs: " & " flag1_187 = "& Convert_SLV_To_Hex_String(flag1_187) & " type_cast_265_wire = "& Convert_SLV_To_Hex_String(type_cast_265_wire) & " konst_266_wire_constant = "& Convert_SLV_To_Hex_String(konst_266_wire_constant) & " outputs:" & " n_word_start_268= "  & Convert_SLV_To_Hex_String(n_word_start_268));
      --
    end process; 
    -- flow-through select operator MUX_267_inst
    n_word_start_268 <= type_cast_265_wire when (flag1_187(0) /=  '0') else konst_266_wire_constant;
    -- logger for split-operator MUX_278_inst flow-through 
    process(n_address_279) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUX_278_inst:flowthrough inputs: " & " flag1_187 = "& Convert_SLV_To_Hex_String(flag1_187) & " type_cast_274_wire = "& Convert_SLV_To_Hex_String(type_cast_274_wire) & " ADD_u64_u64_277_wire = "& Convert_SLV_To_Hex_String(ADD_u64_u64_277_wire) & " outputs:" & " n_address_279= "  & Convert_SLV_To_Hex_String(n_address_279));
      --
    end process; 
    -- flow-through select operator MUX_278_inst
    n_address_279 <= type_cast_274_wire when (flag1_187(0) /=  '0') else ADD_u64_u64_277_wire;
    -- logger for split-operator MUX_286_inst flow-through 
    process(n_left_287) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUX_286_inst:flowthrough inputs: " & " flag1_187 = "& Convert_SLV_To_Hex_String(flag1_187) & " nl_start_34 = "& Convert_SLV_To_Hex_String(nl_start_34) & " SUB_u16_u16_285_wire = "& Convert_SLV_To_Hex_String(SUB_u16_u16_285_wire) & " outputs:" & " n_left_287= "  & Convert_SLV_To_Hex_String(n_left_287));
      --
    end process; 
    -- flow-through select operator MUX_286_inst
    n_left_287 <= nl_start_34 when (flag1_187(0) /=  '0') else SUB_u16_u16_285_wire;
    -- logger for split-operator MUX_299_inst flow-through 
    process(MUX_299_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUX_299_inst:flowthrough inputs: " & " UGT_u16_u1_294_wire = "& Convert_SLV_To_Hex_String(UGT_u16_u1_294_wire) & " SUB_u16_u16_297_wire = "& Convert_SLV_To_Hex_String(SUB_u16_u16_297_wire) & " fn_blk_42 = "& Convert_SLV_To_Hex_String(fn_blk_42) & " outputs:" & " MUX_299_wire= "  & Convert_SLV_To_Hex_String(MUX_299_wire));
      --
    end process; 
    -- flow-through select operator MUX_299_inst
    MUX_299_wire <= SUB_u16_u16_297_wire when (UGT_u16_u1_294_wire(0) /=  '0') else fn_blk_42;
    -- logger for split-operator MUX_305_inst flow-through 
    process(MUX_305_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUX_305_inst:flowthrough inputs: " & " ULT_u16_u1_302_wire = "& Convert_SLV_To_Hex_String(ULT_u16_u1_302_wire) & " n_left_287 = "& Convert_SLV_To_Hex_String(n_left_287) & " konst_304_wire_constant = "& Convert_SLV_To_Hex_String(konst_304_wire_constant) & " outputs:" & " MUX_305_wire= "  & Convert_SLV_To_Hex_String(MUX_305_wire));
      --
    end process; 
    -- flow-through select operator MUX_305_inst
    MUX_305_wire <= n_left_287 when (ULT_u16_u1_302_wire(0) /=  '0') else konst_304_wire_constant;
    -- logger for split-operator MUX_306_inst flow-through 
    process(n_blk_307) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUX_306_inst:flowthrough inputs: " & " flag1_187 = "& Convert_SLV_To_Hex_String(flag1_187) & " MUX_299_wire = "& Convert_SLV_To_Hex_String(MUX_299_wire) & " MUX_305_wire = "& Convert_SLV_To_Hex_String(MUX_305_wire) & " outputs:" & " n_blk_307= "  & Convert_SLV_To_Hex_String(n_blk_307));
      --
    end process; 
    -- flow-through select operator MUX_306_inst
    n_blk_307 <= MUX_299_wire when (flag1_187(0) /=  '0') else MUX_305_wire;
    -- logger for split-operator MUX_41_inst flow-through 
    process(fn_blk_42) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUX_41_inst:flowthrough inputs: " & " ULT_u16_u1_38_wire = "& Convert_SLV_To_Hex_String(ULT_u16_u1_38_wire) & " num_cont_buffer = "& Convert_SLV_To_Hex_String(num_cont_buffer) & " konst_40_wire_constant = "& Convert_SLV_To_Hex_String(konst_40_wire_constant) & " outputs:" & " fn_blk_42= "  & Convert_SLV_To_Hex_String(fn_blk_42));
      --
    end process; 
    -- flow-through select operator MUX_41_inst
    fn_blk_42 <= num_cont_buffer when (ULT_u16_u1_38_wire(0) /=  '0') else konst_40_wire_constant;
    -- logger for split-operator slice_141_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_141_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:slice_141_inst:started:   inputs: " & " word_read_138 = "& Convert_SLV_To_Hex_String(word_read_138));
          --
        end if; 
        if slice_141_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:slice_141_inst:finished:  outputs: " & " w1_142= "  & Convert_SLV_To_Hex_String(w1_142));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_141_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_141_inst_req_0;
      slice_141_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_141_inst_req_1;
      slice_141_inst_ack_1<= update_ack(0);
      slice_141_inst: SliceSplitProtocol generic map(name => "slice_141_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_138, dout => w1_142, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_145_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_145_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:slice_145_inst:started:   inputs: " & " word_read_138 = "& Convert_SLV_To_Hex_String(word_read_138));
          --
        end if; 
        if slice_145_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:slice_145_inst:finished:  outputs: " & " w2_146= "  & Convert_SLV_To_Hex_String(w2_146));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_145_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_145_inst_req_0;
      slice_145_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_145_inst_req_1;
      slice_145_inst_ack_1<= update_ack(0);
      slice_145_inst: SliceSplitProtocol generic map(name => "slice_145_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_138, dout => w2_146, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_149_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_149_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:slice_149_inst:started:   inputs: " & " word_read_138 = "& Convert_SLV_To_Hex_String(word_read_138));
          --
        end if; 
        if slice_149_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:slice_149_inst:finished:  outputs: " & " w3_150= "  & Convert_SLV_To_Hex_String(w3_150));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_149_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_149_inst_req_0;
      slice_149_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_149_inst_req_1;
      slice_149_inst_ack_1<= update_ack(0);
      slice_149_inst: SliceSplitProtocol generic map(name => "slice_149_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_138, dout => w3_150, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_153_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_153_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:slice_153_inst:started:   inputs: " & " word_read_138 = "& Convert_SLV_To_Hex_String(word_read_138));
          --
        end if; 
        if slice_153_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:slice_153_inst:finished:  outputs: " & " w4_154= "  & Convert_SLV_To_Hex_String(w4_154));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_153_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_153_inst_req_0;
      slice_153_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_153_inst_req_1;
      slice_153_inst_ack_1<= update_ack(0);
      slice_153_inst: SliceSplitProtocol generic map(name => "slice_153_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_138, dout => w4_154, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator W_c1_155_delayed_14_0_155_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_c1_155_delayed_14_0_155_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:W_c1_155_delayed_14_0_155_inst:started:   inputs: " & " c1_85 = "& Convert_SLV_To_Hex_String(c1_85));
          --
        end if; 
        if W_c1_155_delayed_14_0_155_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:W_c1_155_delayed_14_0_155_inst:finished:  outputs: " & " c1_155_delayed_14_0_157= "  & Convert_SLV_To_Hex_String(c1_155_delayed_14_0_157));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_c1_155_delayed_14_0_155_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c1_155_delayed_14_0_155_inst_req_0;
      W_c1_155_delayed_14_0_155_inst_ack_0<= wack(0);
      rreq(0) <= W_c1_155_delayed_14_0_155_inst_req_1;
      W_c1_155_delayed_14_0_155_inst_ack_1<= rack(0);
      W_c1_155_delayed_14_0_155_inst : InterlockBuffer generic map ( -- 
        name => "W_c1_155_delayed_14_0_155_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c1_85,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c1_155_delayed_14_0_157,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_c2_159_delayed_14_0_162_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_c2_159_delayed_14_0_162_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:W_c2_159_delayed_14_0_162_inst:started:   inputs: " & " c2_98 = "& Convert_SLV_To_Hex_String(c2_98));
          --
        end if; 
        if W_c2_159_delayed_14_0_162_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:W_c2_159_delayed_14_0_162_inst:finished:  outputs: " & " c2_159_delayed_14_0_164= "  & Convert_SLV_To_Hex_String(c2_159_delayed_14_0_164));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_c2_159_delayed_14_0_162_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c2_159_delayed_14_0_162_inst_req_0;
      W_c2_159_delayed_14_0_162_inst_ack_0<= wack(0);
      rreq(0) <= W_c2_159_delayed_14_0_162_inst_req_1;
      W_c2_159_delayed_14_0_162_inst_ack_1<= rack(0);
      W_c2_159_delayed_14_0_162_inst : InterlockBuffer generic map ( -- 
        name => "W_c2_159_delayed_14_0_162_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c2_98,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c2_159_delayed_14_0_164,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_c3_163_delayed_14_0_169_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_c3_163_delayed_14_0_169_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:W_c3_163_delayed_14_0_169_inst:started:   inputs: " & " c3_119 = "& Convert_SLV_To_Hex_String(c3_119));
          --
        end if; 
        if W_c3_163_delayed_14_0_169_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:W_c3_163_delayed_14_0_169_inst:finished:  outputs: " & " c3_163_delayed_14_0_171= "  & Convert_SLV_To_Hex_String(c3_163_delayed_14_0_171));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_c3_163_delayed_14_0_169_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c3_163_delayed_14_0_169_inst_req_0;
      W_c3_163_delayed_14_0_169_inst_ack_0<= wack(0);
      rreq(0) <= W_c3_163_delayed_14_0_169_inst_req_1;
      W_c3_163_delayed_14_0_169_inst_ack_1<= rack(0);
      W_c3_163_delayed_14_0_169_inst : InterlockBuffer generic map ( -- 
        name => "W_c3_163_delayed_14_0_169_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c3_119,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c3_163_delayed_14_0_171,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_c4_167_delayed_14_0_176_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_c4_167_delayed_14_0_176_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:W_c4_167_delayed_14_0_176_inst:started:   inputs: " & " c4_127 = "& Convert_SLV_To_Hex_String(c4_127));
          --
        end if; 
        if W_c4_167_delayed_14_0_176_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:W_c4_167_delayed_14_0_176_inst:finished:  outputs: " & " c4_167_delayed_14_0_178= "  & Convert_SLV_To_Hex_String(c4_167_delayed_14_0_178));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_c4_167_delayed_14_0_176_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c4_167_delayed_14_0_176_inst_req_0;
      W_c4_167_delayed_14_0_176_inst_ack_0<= wack(0);
      rreq(0) <= W_c4_167_delayed_14_0_176_inst_req_1;
      W_c4_167_delayed_14_0_176_inst_ack_1<= rack(0);
      W_c4_167_delayed_14_0_176_inst : InterlockBuffer generic map ( -- 
        name => "W_c4_167_delayed_14_0_176_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c4_127,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c4_167_delayed_14_0_178,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_nl_start_32_inst flow-through 
    process(nl_start_34) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:W_nl_start_32_inst:flowthrough inputs: " & " num_cont_buffer = "& Convert_SLV_To_Hex_String(num_cont_buffer) & " outputs:" & " nl_start_34= "  & Convert_SLV_To_Hex_String(nl_start_34));
      --
    end process; 
    -- interlock W_nl_start_32_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := num_cont_buffer(15 downto 0);
      nl_start_34 <= tmp_var; -- 
    end process;
    -- logger for split-operator addr_of_133_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_133_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:addr_of_133_final_reg:started:   inputs: " & " array_obj_ref_132_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_132_root_address));
          --
        end if; 
        if addr_of_133_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:addr_of_133_final_reg:finished:  outputs: " & " fetch_addr_134= "  & Convert_SLV_To_Hex_String(fetch_addr_134));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_133_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_133_final_reg_req_0;
      addr_of_133_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_133_final_reg_req_1;
      addr_of_133_final_reg_ack_1<= rack(0);
      addr_of_133_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_133_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_132_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_134,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_address_279_47_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_address_279_47_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_address_279_47_buf:started:   inputs: " & " n_address_279 = "& Convert_SLV_To_Hex_String(n_address_279));
          --
        end if; 
        if n_address_279_47_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_address_279_47_buf:finished:  outputs: " & " n_address_279_47_buffered= "  & Convert_SLV_To_Hex_String(n_address_279_47_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_address_279_47_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address_279_47_buf_req_0;
      n_address_279_47_buf_ack_0<= wack(0);
      rreq(0) <= n_address_279_47_buf_req_1;
      n_address_279_47_buf_ack_1<= rack(0);
      n_address_279_47_buf : InterlockBuffer generic map ( -- 
        name => "n_address_279_47_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address_279,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address_279_47_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_blk_307_62_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_blk_307_62_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_blk_307_62_buf:started:   inputs: " & " n_blk_307 = "& Convert_SLV_To_Hex_String(n_blk_307));
          --
        end if; 
        if n_blk_307_62_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_blk_307_62_buf:finished:  outputs: " & " n_blk_307_62_buffered= "  & Convert_SLV_To_Hex_String(n_blk_307_62_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_blk_307_62_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_blk_307_62_buf_req_0;
      n_blk_307_62_buf_ack_0<= wack(0);
      rreq(0) <= n_blk_307_62_buf_req_1;
      n_blk_307_62_buf_ack_1<= rack(0);
      n_blk_307_62_buf : InterlockBuffer generic map ( -- 
        name => "n_blk_307_62_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_blk_307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_blk_307_62_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_col_221_74_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_col_221_74_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_col_221_74_buf:started:   inputs: " & " n_col_221 = "& Convert_SLV_To_Hex_String(n_col_221));
          --
        end if; 
        if n_col_221_74_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_col_221_74_buf:finished:  outputs: " & " n_col_221_74_buffered= "  & Convert_SLV_To_Hex_String(n_col_221_74_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_col_221_74_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_221_74_buf_req_0;
      n_col_221_74_buf_ack_0<= wack(0);
      rreq(0) <= n_col_221_74_buf_req_1;
      n_col_221_74_buf_ack_1<= rack(0);
      n_col_221_74_buf : InterlockBuffer generic map ( -- 
        name => "n_col_221_74_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_221,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_221_74_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_left_287_59_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_left_287_59_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_left_287_59_buf:started:   inputs: " & " n_left_287 = "& Convert_SLV_To_Hex_String(n_left_287));
          --
        end if; 
        if n_left_287_59_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_left_287_59_buf:finished:  outputs: " & " n_left_287_59_buffered= "  & Convert_SLV_To_Hex_String(n_left_287_59_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_left_287_59_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_left_287_59_buf_req_0;
      n_left_287_59_buf_ack_0<= wack(0);
      rreq(0) <= n_left_287_59_buf_req_1;
      n_left_287_59_buf_ack_1<= rack(0);
      n_left_287_59_buf : InterlockBuffer generic map ( -- 
        name => "n_left_287_59_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_left_287,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_left_287_59_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_row_233_77_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_row_233_77_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_row_233_77_buf:started:   inputs: " & " n_row_233 = "& Convert_SLV_To_Hex_String(n_row_233));
          --
        end if; 
        if n_row_233_77_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_row_233_77_buf:finished:  outputs: " & " n_row_233_77_buffered= "  & Convert_SLV_To_Hex_String(n_row_233_77_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_row_233_77_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_233_77_buf_req_0;
      n_row_233_77_buf_ack_0<= wack(0);
      rreq(0) <= n_row_233_77_buf_req_1;
      n_row_233_77_buf_ack_1<= rack(0);
      n_row_233_77_buf : InterlockBuffer generic map ( -- 
        name => "n_row_233_77_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_233,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_233_77_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_winr_208_69_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_winr_208_69_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_winr_208_69_buf:started:   inputs: " & " n_winr_208 = "& Convert_SLV_To_Hex_String(n_winr_208));
          --
        end if; 
        if n_winr_208_69_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_winr_208_69_buf:finished:  outputs: " & " n_winr_208_69_buffered= "  & Convert_SLV_To_Hex_String(n_winr_208_69_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_winr_208_69_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_winr_208_69_buf_req_0;
      n_winr_208_69_buf_ack_0<= wack(0);
      rreq(0) <= n_winr_208_69_buf_req_1;
      n_winr_208_69_buf_ack_1<= rack(0);
      n_winr_208_69_buf : InterlockBuffer generic map ( -- 
        name => "n_winr_208_69_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_winr_208,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_winr_208_69_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_word_start_268_52_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_word_start_268_52_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_word_start_268_52_buf:started:   inputs: " & " n_word_start_268 = "& Convert_SLV_To_Hex_String(n_word_start_268));
          --
        end if; 
        if n_word_start_268_52_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:n_word_start_268_52_buf:finished:  outputs: " & " n_word_start_268_52_buffered= "  & Convert_SLV_To_Hex_String(n_word_start_268_52_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_word_start_268_52_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_word_start_268_52_buf_req_0;
      n_word_start_268_52_buf_ack_0<= wack(0);
      rreq(0) <= n_word_start_268_52_buf_req_1;
      n_word_start_268_52_buf_ack_1<= rack(0);
      n_word_start_268_52_buf : InterlockBuffer generic map ( -- 
        name => "n_word_start_268_52_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_word_start_268,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_word_start_268_52_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator nl_start_34_58_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if nl_start_34_58_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:nl_start_34_58_buf:started:   inputs: " & " nl_start_34 = "& Convert_SLV_To_Hex_String(nl_start_34));
          --
        end if; 
        if nl_start_34_58_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:nl_start_34_58_buf:finished:  outputs: " & " nl_start_34_58_buffered= "  & Convert_SLV_To_Hex_String(nl_start_34_58_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    nl_start_34_58_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nl_start_34_58_buf_req_0;
      nl_start_34_58_buf_ack_0<= wack(0);
      rreq(0) <= nl_start_34_58_buf_req_1;
      nl_start_34_58_buf_ack_1<= rack(0);
      nl_start_34_58_buf : InterlockBuffer generic map ( -- 
        name => "nl_start_34_58_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nl_start_34,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nl_start_34_58_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_123_inst flow-through 
    process(type_cast_123_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:type_cast_123_inst:flowthrough inputs: " & " word_start_50 = "& Convert_SLV_To_Hex_String(word_start_50) & " outputs:" & " type_cast_123_wire= "  & Convert_SLV_To_Hex_String(type_cast_123_wire));
      --
    end process; 
    -- interlock type_cast_123_inst
    process(word_start_50) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := word_start_50(1 downto 0);
      type_cast_123_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_242_inst flow-through 
    process(na1_243) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:type_cast_242_inst:flowthrough inputs: " & " MUL_u16_u16_241_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_241_wire) & " outputs:" & " na1_243= "  & Convert_SLV_To_Hex_String(na1_243));
      --
    end process; 
    -- interlock type_cast_242_inst
    process(MUL_u16_u16_241_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_241_wire(15 downto 0);
      na1_243 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_247_inst flow-through 
    process(type_cast_247_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:type_cast_247_inst:flowthrough inputs: " & " n_winr_208 = "& Convert_SLV_To_Hex_String(n_winr_208) & " outputs:" & " type_cast_247_wire= "  & Convert_SLV_To_Hex_String(type_cast_247_wire));
      --
    end process; 
    -- interlock type_cast_247_inst
    process(n_winr_208) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_winr_208(15 downto 0);
      type_cast_247_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_249_inst flow-through 
    process(na2_250) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:type_cast_249_inst:flowthrough inputs: " & " MUL_u32_u32_248_wire = "& Convert_SLV_To_Hex_String(MUL_u32_u32_248_wire) & " outputs:" & " na2_250= "  & Convert_SLV_To_Hex_String(na2_250));
      --
    end process; 
    -- interlock type_cast_249_inst
    process(MUL_u32_u32_248_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := MUL_u32_u32_248_wire(31 downto 0);
      na2_250 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_260_inst flow-through 
    process(na4_261) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:type_cast_260_inst:flowthrough inputs: " & " AND_u32_u32_259_wire = "& Convert_SLV_To_Hex_String(AND_u32_u32_259_wire) & " outputs:" & " na4_261= "  & Convert_SLV_To_Hex_String(na4_261));
      --
    end process; 
    -- interlock type_cast_260_inst
    process(AND_u32_u32_259_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := AND_u32_u32_259_wire(15 downto 0);
      na4_261 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_265_inst flow-through 
    process(type_cast_265_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:type_cast_265_inst:flowthrough inputs: " & " na4_261 = "& Convert_SLV_To_Hex_String(na4_261) & " outputs:" & " type_cast_265_wire= "  & Convert_SLV_To_Hex_String(type_cast_265_wire));
      --
    end process; 
    -- interlock type_cast_265_inst
    process(na4_261) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := na4_261(1 downto 0);
      type_cast_265_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_274_inst flow-through 
    process(type_cast_274_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:type_cast_274_inst:flowthrough inputs: " & " LSHR_u32_u32_273_wire = "& Convert_SLV_To_Hex_String(LSHR_u32_u32_273_wire) & " outputs:" & " type_cast_274_wire= "  & Convert_SLV_To_Hex_String(type_cast_274_wire));
      --
    end process; 
    -- interlock type_cast_274_inst
    process(LSHR_u32_u32_273_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_273_wire(31 downto 0);
      type_cast_274_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_30_inst flow-through 
    process(m_factor_31) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:type_cast_30_inst:flowthrough inputs: " & " MUL_u16_u16_29_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_29_wire) & " outputs:" & " m_factor_31= "  & Convert_SLV_To_Hex_String(m_factor_31));
      --
    end process; 
    -- interlock type_cast_30_inst
    process(MUL_u16_u16_29_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_29_wire(15 downto 0);
      m_factor_31 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_64_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_64_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:type_cast_64_inst:started:   inputs: " & " fn_blk_42 = "& Convert_SLV_To_Hex_String(fn_blk_42));
          --
        end if; 
        if type_cast_64_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:type_cast_64_inst:finished:  outputs: " & " type_cast_64_wire= "  & Convert_SLV_To_Hex_String(type_cast_64_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_64_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_64_inst_req_0;
      type_cast_64_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_64_inst_req_1;
      type_cast_64_inst_ack_1<= rack(0);
      type_cast_64_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_64_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_blk_42,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_64_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_132_index_1_rename flow-through 
    process(R_address_131_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:array_obj_ref_132_index_1_rename:flowthrough  inputs: " & " R_address_131_resized = "& Convert_SLV_To_Hex_String(R_address_131_resized) & "outputs: " & " R_address_131_scaled= "  & Convert_SLV_To_Hex_String(R_address_131_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_132_index_1_rename
    process(R_address_131_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_131_resized;
      ov(13 downto 0) := iv;
      R_address_131_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_132_index_1_resize flow-through 
    process(R_address_131_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:array_obj_ref_132_index_1_resize:flowthrough  inputs: " & " address_45 = "& Convert_SLV_To_Hex_String(address_45) & "outputs: " & " R_address_131_resized= "  & Convert_SLV_To_Hex_String(R_address_131_resized));
      --
    end process; 
    -- equivalence array_obj_ref_132_index_1_resize
    process(address_45) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_45;
      ov := iv(13 downto 0);
      R_address_131_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_132_root_address_inst flow-through 
    process(array_obj_ref_132_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:array_obj_ref_132_root_address_inst:flowthrough  inputs: " & " array_obj_ref_132_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_132_final_offset) & "outputs: " & " array_obj_ref_132_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_132_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_132_root_address_inst
    process(array_obj_ref_132_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_132_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_132_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_137_addr_0 flow-through 
    process(ptr_deref_137_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ptr_deref_137_addr_0:flowthrough  inputs: " & " ptr_deref_137_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_137_root_address) & "outputs: " & " ptr_deref_137_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_137_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_137_addr_0
    process(ptr_deref_137_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_137_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_137_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_137_base_resize flow-through 
    process(ptr_deref_137_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ptr_deref_137_base_resize:flowthrough  inputs: " & " fetch_addr_134 = "& Convert_SLV_To_Hex_String(fetch_addr_134) & "outputs: " & " ptr_deref_137_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_137_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_137_base_resize
    process(fetch_addr_134) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_134;
      ov := iv(13 downto 0);
      ptr_deref_137_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_137_gather_scatter flow-through 
    process(word_read_138) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ptr_deref_137_gather_scatter:flowthrough  inputs: " & " ptr_deref_137_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_137_data_0) & "outputs: " & " word_read_138= "  & Convert_SLV_To_Hex_String(word_read_138));
      --
    end process; 
    -- equivalence ptr_deref_137_gather_scatter
    process(ptr_deref_137_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_137_data_0;
      ov(63 downto 0) := iv;
      word_read_138 <= ov(63 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_137_root_address_inst flow-through 
    process(ptr_deref_137_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ptr_deref_137_root_address_inst:flowthrough  inputs: " & " ptr_deref_137_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_137_resized_base_address) & "outputs: " & " ptr_deref_137_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_137_root_address));
      --
    end process; 
    -- equivalence ptr_deref_137_root_address_inst
    process(ptr_deref_137_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_137_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_137_root_address <= ov(13 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_43_branch_req_0," req0 do_while_stmt_43_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_43_branch_ack_0," ack0 do_while_stmt_43_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_43_branch_ack_1," ack1 do_while_stmt_43_branch");
    do_while_stmt_43_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NEQ_u16_u1_311_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_43_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_43_branch_req_0,
          ack0 => do_while_stmt_43_branch_ack_0,
          ack1 => do_while_stmt_43_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u16_u16_124_inst flow-through 
    process(ADD_u16_u16_124_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ADD_u16_u16_124_inst:flowthrough inputs: " & " num_blk_60 = "& Convert_SLV_To_Hex_String(num_blk_60) & " type_cast_123_wire = "& Convert_SLV_To_Hex_String(type_cast_123_wire) & " outputs:" & " ADD_u16_u16_124_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_124_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_124_inst
    process(num_blk_60, type_cast_123_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_blk_60, type_cast_123_wire, tmp_var);
      ADD_u16_u16_124_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_204_inst flow-through 
    process(ADD_u16_u16_204_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ADD_u16_u16_204_inst:flowthrough inputs: " & " winr_65 = "& Convert_SLV_To_Hex_String(winr_65) & " konst_203_wire_constant = "& Convert_SLV_To_Hex_String(konst_203_wire_constant) & " outputs:" & " ADD_u16_u16_204_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_204_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_204_inst
    process(winr_65) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(winr_65, konst_203_wire_constant, tmp_var);
      ADD_u16_u16_204_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_217_inst flow-through 
    process(ADD_u16_u16_217_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ADD_u16_u16_217_inst:flowthrough inputs: " & " col_70 = "& Convert_SLV_To_Hex_String(col_70) & " konst_216_wire_constant = "& Convert_SLV_To_Hex_String(konst_216_wire_constant) & " outputs:" & " ADD_u16_u16_217_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_217_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_217_inst
    process(col_70) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_70, konst_216_wire_constant, tmp_var);
      ADD_u16_u16_217_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_230_inst flow-through 
    process(ADD_u16_u16_230_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ADD_u16_u16_230_inst:flowthrough inputs: " & " row_75 = "& Convert_SLV_To_Hex_String(row_75) & " konst_229_wire_constant = "& Convert_SLV_To_Hex_String(konst_229_wire_constant) & " outputs:" & " ADD_u16_u16_230_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_230_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_230_inst
    process(row_75) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_75, konst_229_wire_constant, tmp_var);
      ADD_u16_u16_230_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_240_inst flow-through 
    process(ADD_u16_u16_240_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ADD_u16_u16_240_inst:flowthrough inputs: " & " n_col_221 = "& Convert_SLV_To_Hex_String(n_col_221) & " MUL_u16_u16_239_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_239_wire) & " outputs:" & " ADD_u16_u16_240_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_240_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_240_inst
    process(n_col_221, MUL_u16_u16_239_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(n_col_221, MUL_u16_u16_239_wire, tmp_var);
      ADD_u16_u16_240_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_292_inst flow-through 
    process(ADD_u16_u16_292_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ADD_u16_u16_292_inst:flowthrough inputs: " & " fn_blk_42 = "& Convert_SLV_To_Hex_String(fn_blk_42) & " na4_261 = "& Convert_SLV_To_Hex_String(na4_261) & " outputs:" & " ADD_u16_u16_292_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_292_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_292_inst
    process(fn_blk_42, na4_261) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(fn_blk_42, na4_261, tmp_var);
      ADD_u16_u16_292_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_254_inst flow-through 
    process(na3_255) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ADD_u32_u32_254_inst:flowthrough inputs: " & " na1_243 = "& Convert_SLV_To_Hex_String(na1_243) & " na2_250 = "& Convert_SLV_To_Hex_String(na2_250) & " outputs:" & " na3_255= "  & Convert_SLV_To_Hex_String(na3_255));
      --
    end process; 
    -- binary operator ADD_u32_u32_254_inst
    process(na1_243, na2_250) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(na1_243, na2_250, tmp_var);
      na3_255 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u64_u64_277_inst flow-through 
    process(ADD_u64_u64_277_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ADD_u64_u64_277_inst:flowthrough inputs: " & " address_45 = "& Convert_SLV_To_Hex_String(address_45) & " konst_276_wire_constant = "& Convert_SLV_To_Hex_String(konst_276_wire_constant) & " outputs:" & " ADD_u64_u64_277_wire= "  & Convert_SLV_To_Hex_String(ADD_u64_u64_277_wire));
      --
    end process; 
    -- binary operator ADD_u64_u64_277_inst
    process(address_45) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address_45, konst_276_wire_constant, tmp_var);
      ADD_u64_u64_277_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_106_inst flow-through 
    process(AND_u1_u1_106_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:AND_u1_u1_106_inst:flowthrough inputs: " & " EQ_u2_u1_102_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_102_wire) & " UGT_u16_u1_105_wire = "& Convert_SLV_To_Hex_String(UGT_u16_u1_105_wire) & " outputs:" & " AND_u1_u1_106_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_106_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_106_inst
    process(EQ_u2_u1_102_wire, UGT_u16_u1_105_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_102_wire, UGT_u16_u1_105_wire, tmp_var);
      AND_u1_u1_106_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_113_inst flow-through 
    process(AND_u1_u1_113_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:AND_u1_u1_113_inst:flowthrough inputs: " & " EQ_u2_u1_109_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_109_wire) & " UGT_u16_u1_112_wire = "& Convert_SLV_To_Hex_String(UGT_u16_u1_112_wire) & " outputs:" & " AND_u1_u1_113_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_113_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_113_inst
    process(EQ_u2_u1_109_wire, UGT_u16_u1_112_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_109_wire, UGT_u16_u1_112_wire, tmp_var);
      AND_u1_u1_113_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_212_inst flow-through 
    process(AND_u1_u1_212_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:AND_u1_u1_212_inst:flowthrough inputs: " & " winr_done_192 = "& Convert_SLV_To_Hex_String(winr_done_192) & " flag1_187 = "& Convert_SLV_To_Hex_String(flag1_187) & " outputs:" & " AND_u1_u1_212_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_212_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_212_inst
    process(winr_done_192, flag1_187) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_192, flag1_187, tmp_var);
      AND_u1_u1_212_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_226_inst flow-through 
    process(AND_u1_u1_226_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:AND_u1_u1_226_inst:flowthrough inputs: " & " col_done_197 = "& Convert_SLV_To_Hex_String(col_done_197) & " flag1_187 = "& Convert_SLV_To_Hex_String(flag1_187) & " outputs:" & " AND_u1_u1_226_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_226_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_226_inst
    process(col_done_197, flag1_187) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_197, flag1_187, tmp_var);
      AND_u1_u1_226_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_227_inst flow-through 
    process(AND_u1_u1_227_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:AND_u1_u1_227_inst:flowthrough inputs: " & " winr_done_192 = "& Convert_SLV_To_Hex_String(winr_done_192) & " AND_u1_u1_226_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_226_wire) & " outputs:" & " AND_u1_u1_227_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_227_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_227_inst
    process(winr_done_192, AND_u1_u1_226_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_192, AND_u1_u1_226_wire, tmp_var);
      AND_u1_u1_227_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_93_inst flow-through 
    process(AND_u1_u1_93_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:AND_u1_u1_93_inst:flowthrough inputs: " & " EQ_u2_u1_89_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_89_wire) & " UGT_u16_u1_92_wire = "& Convert_SLV_To_Hex_String(UGT_u16_u1_92_wire) & " outputs:" & " AND_u1_u1_93_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_93_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_93_inst
    process(EQ_u2_u1_89_wire, UGT_u16_u1_92_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_89_wire, UGT_u16_u1_92_wire, tmp_var);
      AND_u1_u1_93_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u32_u32_259_inst flow-through 
    process(AND_u32_u32_259_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:AND_u32_u32_259_inst:flowthrough inputs: " & " na3_255 = "& Convert_SLV_To_Hex_String(na3_255) & " konst_258_wire_constant = "& Convert_SLV_To_Hex_String(konst_258_wire_constant) & " outputs:" & " AND_u32_u32_259_wire= "  & Convert_SLV_To_Hex_String(AND_u32_u32_259_wire));
      --
    end process; 
    -- binary operator AND_u32_u32_259_inst
    process(na3_255) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(na3_255, konst_258_wire_constant, tmp_var);
      AND_u32_u32_259_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u16_u1_186_inst flow-through 
    process(flag1_187) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:EQ_u16_u1_186_inst:flowthrough inputs: " & " num_left_56 = "& Convert_SLV_To_Hex_String(num_left_56) & " num_blk_60 = "& Convert_SLV_To_Hex_String(num_blk_60) & " outputs:" & " flag1_187= "  & Convert_SLV_To_Hex_String(flag1_187));
      --
    end process; 
    -- binary operator EQ_u16_u1_186_inst
    process(num_left_56, num_blk_60) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_left_56, num_blk_60, tmp_var);
      flag1_187 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u16_u1_191_inst flow-through 
    process(winr_done_192) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:EQ_u16_u1_191_inst:flowthrough inputs: " & " winr_65 = "& Convert_SLV_To_Hex_String(winr_65) & " rk1_buffer = "& Convert_SLV_To_Hex_String(rk1_buffer) & " outputs:" & " winr_done_192= "  & Convert_SLV_To_Hex_String(winr_done_192));
      --
    end process; 
    -- binary operator EQ_u16_u1_191_inst
    process(winr_65, rk1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(winr_65, rk1_buffer, tmp_var);
      winr_done_192 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u16_u1_196_inst flow-through 
    process(col_done_197) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:EQ_u16_u1_196_inst:flowthrough inputs: " & " col_70 = "& Convert_SLV_To_Hex_String(col_70) & " col1_buffer = "& Convert_SLV_To_Hex_String(col1_buffer) & " outputs:" & " col_done_197= "  & Convert_SLV_To_Hex_String(col_done_197));
      --
    end process; 
    -- binary operator EQ_u16_u1_196_inst
    process(col_70, col1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_70, col1_buffer, tmp_var);
      col_done_197 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_102_inst flow-through 
    process(EQ_u2_u1_102_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:EQ_u2_u1_102_inst:flowthrough inputs: " & " word_start_50 = "& Convert_SLV_To_Hex_String(word_start_50) & " konst_101_wire_constant = "& Convert_SLV_To_Hex_String(konst_101_wire_constant) & " outputs:" & " EQ_u2_u1_102_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_102_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_102_inst
    process(word_start_50) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_50, konst_101_wire_constant, tmp_var);
      EQ_u2_u1_102_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_109_inst flow-through 
    process(EQ_u2_u1_109_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:EQ_u2_u1_109_inst:flowthrough inputs: " & " word_start_50 = "& Convert_SLV_To_Hex_String(word_start_50) & " konst_108_wire_constant = "& Convert_SLV_To_Hex_String(konst_108_wire_constant) & " outputs:" & " EQ_u2_u1_109_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_109_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_109_inst
    process(word_start_50) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_50, konst_108_wire_constant, tmp_var);
      EQ_u2_u1_109_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_116_inst flow-through 
    process(EQ_u2_u1_116_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:EQ_u2_u1_116_inst:flowthrough inputs: " & " word_start_50 = "& Convert_SLV_To_Hex_String(word_start_50) & " konst_115_wire_constant = "& Convert_SLV_To_Hex_String(konst_115_wire_constant) & " outputs:" & " EQ_u2_u1_116_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_116_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_116_inst
    process(word_start_50) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_50, konst_115_wire_constant, tmp_var);
      EQ_u2_u1_116_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_84_inst flow-through 
    process(c1_85) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:EQ_u2_u1_84_inst:flowthrough inputs: " & " word_start_50 = "& Convert_SLV_To_Hex_String(word_start_50) & " konst_83_wire_constant = "& Convert_SLV_To_Hex_String(konst_83_wire_constant) & " outputs:" & " c1_85= "  & Convert_SLV_To_Hex_String(c1_85));
      --
    end process; 
    -- binary operator EQ_u2_u1_84_inst
    process(word_start_50) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_50, konst_83_wire_constant, tmp_var);
      c1_85 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_89_inst flow-through 
    process(EQ_u2_u1_89_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:EQ_u2_u1_89_inst:flowthrough inputs: " & " word_start_50 = "& Convert_SLV_To_Hex_String(word_start_50) & " konst_88_wire_constant = "& Convert_SLV_To_Hex_String(konst_88_wire_constant) & " outputs:" & " EQ_u2_u1_89_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_89_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_89_inst
    process(word_start_50) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_50, konst_88_wire_constant, tmp_var);
      EQ_u2_u1_89_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_96_inst flow-through 
    process(EQ_u2_u1_96_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:EQ_u2_u1_96_inst:flowthrough inputs: " & " word_start_50 = "& Convert_SLV_To_Hex_String(word_start_50) & " konst_95_wire_constant = "& Convert_SLV_To_Hex_String(konst_95_wire_constant) & " outputs:" & " EQ_u2_u1_96_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_96_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_96_inst
    process(word_start_50) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_50, konst_95_wire_constant, tmp_var);
      EQ_u2_u1_96_wire <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u32_u32_273_inst flow-through 
    process(LSHR_u32_u32_273_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:LSHR_u32_u32_273_inst:flowthrough inputs: " & " na3_255 = "& Convert_SLV_To_Hex_String(na3_255) & " konst_272_wire_constant = "& Convert_SLV_To_Hex_String(konst_272_wire_constant) & " outputs:" & " LSHR_u32_u32_273_wire= "  & Convert_SLV_To_Hex_String(LSHR_u32_u32_273_wire));
      --
    end process; 
    -- binary operator LSHR_u32_u32_273_inst
    process(na3_255) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(na3_255, konst_272_wire_constant, tmp_var);
      LSHR_u32_u32_273_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_239_inst flow-through 
    process(MUL_u16_u16_239_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUL_u16_u16_239_inst:flowthrough inputs: " & " ct_buffer = "& Convert_SLV_To_Hex_String(ct_buffer) & " n_row_233 = "& Convert_SLV_To_Hex_String(n_row_233) & " outputs:" & " MUL_u16_u16_239_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_239_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_239_inst
    process(ct_buffer, n_row_233) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, n_row_233, tmp_var);
      MUL_u16_u16_239_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_241_inst flow-through 
    process(MUL_u16_u16_241_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUL_u16_u16_241_inst:flowthrough inputs: " & " chl_in_buffer = "& Convert_SLV_To_Hex_String(chl_in_buffer) & " ADD_u16_u16_240_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_240_wire) & " outputs:" & " MUL_u16_u16_241_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_241_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_241_inst
    process(chl_in_buffer, ADD_u16_u16_240_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(chl_in_buffer, ADD_u16_u16_240_wire, tmp_var);
      MUL_u16_u16_241_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_29_inst flow-through 
    process(MUL_u16_u16_29_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUL_u16_u16_29_inst:flowthrough inputs: " & " ct_buffer = "& Convert_SLV_To_Hex_String(ct_buffer) & " chl_in_buffer = "& Convert_SLV_To_Hex_String(chl_in_buffer) & " outputs:" & " MUL_u16_u16_29_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_29_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_29_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_29_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u32_u32_248_inst flow-through 
    process(MUL_u32_u32_248_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:MUL_u32_u32_248_inst:flowthrough inputs: " & " m_factor_31 = "& Convert_SLV_To_Hex_String(m_factor_31) & " type_cast_247_wire = "& Convert_SLV_To_Hex_String(type_cast_247_wire) & " outputs:" & " MUL_u32_u32_248_wire= "  & Convert_SLV_To_Hex_String(MUL_u32_u32_248_wire));
      --
    end process; 
    -- binary operator MUL_u32_u32_248_inst
    process(m_factor_31, type_cast_247_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(m_factor_31, type_cast_247_wire, tmp_var);
      MUL_u32_u32_248_wire <= tmp_var; --
    end process;
    -- logger for split-operator NEQ_u16_u1_311_inst flow-through 
    process(NEQ_u16_u1_311_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:NEQ_u16_u1_311_inst:flowthrough inputs: " & " n_row_233 = "& Convert_SLV_To_Hex_String(n_row_233) & " row1_buffer = "& Convert_SLV_To_Hex_String(row1_buffer) & " outputs:" & " NEQ_u16_u1_311_wire= "  & Convert_SLV_To_Hex_String(NEQ_u16_u1_311_wire));
      --
    end process; 
    -- binary operator NEQ_u16_u1_311_inst
    process(n_row_233, row1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(n_row_233, row1_buffer, tmp_var);
      NEQ_u16_u1_311_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_117_inst flow-through 
    process(OR_u1_u1_117_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:OR_u1_u1_117_inst:flowthrough inputs: " & " AND_u1_u1_113_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_113_wire) & " EQ_u2_u1_116_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_116_wire) & " outputs:" & " OR_u1_u1_117_wire= "  & Convert_SLV_To_Hex_String(OR_u1_u1_117_wire));
      --
    end process; 
    -- binary operator OR_u1_u1_117_inst
    process(AND_u1_u1_113_wire, EQ_u2_u1_116_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_113_wire, EQ_u2_u1_116_wire, tmp_var);
      OR_u1_u1_117_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_118_inst flow-through 
    process(c3_119) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:OR_u1_u1_118_inst:flowthrough inputs: " & " AND_u1_u1_106_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_106_wire) & " OR_u1_u1_117_wire = "& Convert_SLV_To_Hex_String(OR_u1_u1_117_wire) & " outputs:" & " c3_119= "  & Convert_SLV_To_Hex_String(c3_119));
      --
    end process; 
    -- binary operator OR_u1_u1_118_inst
    process(AND_u1_u1_106_wire, OR_u1_u1_117_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_106_wire, OR_u1_u1_117_wire, tmp_var);
      c3_119 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_97_inst flow-through 
    process(c2_98) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:OR_u1_u1_97_inst:flowthrough inputs: " & " AND_u1_u1_93_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_93_wire) & " EQ_u2_u1_96_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_96_wire) & " outputs:" & " c2_98= "  & Convert_SLV_To_Hex_String(c2_98));
      --
    end process; 
    -- binary operator OR_u1_u1_97_inst
    process(AND_u1_u1_93_wire, EQ_u2_u1_96_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_93_wire, EQ_u2_u1_96_wire, tmp_var);
      c2_98 <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u16_u16_285_inst flow-through 
    process(SUB_u16_u16_285_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:SUB_u16_u16_285_inst:flowthrough inputs: " & " num_left_56 = "& Convert_SLV_To_Hex_String(num_left_56) & " num_blk_60 = "& Convert_SLV_To_Hex_String(num_blk_60) & " outputs:" & " SUB_u16_u16_285_wire= "  & Convert_SLV_To_Hex_String(SUB_u16_u16_285_wire));
      --
    end process; 
    -- binary operator SUB_u16_u16_285_inst
    process(num_left_56, num_blk_60) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(num_left_56, num_blk_60, tmp_var);
      SUB_u16_u16_285_wire <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u16_u16_297_inst flow-through 
    process(SUB_u16_u16_297_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:SUB_u16_u16_297_inst:flowthrough inputs: " & " konst_295_wire_constant = "& Convert_SLV_To_Hex_String(konst_295_wire_constant) & " na4_261 = "& Convert_SLV_To_Hex_String(na4_261) & " outputs:" & " SUB_u16_u16_297_wire= "  & Convert_SLV_To_Hex_String(SUB_u16_u16_297_wire));
      --
    end process; 
    -- binary operator SUB_u16_u16_297_inst
    process(konst_295_wire_constant, na4_261) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_295_wire_constant, na4_261, tmp_var);
      SUB_u16_u16_297_wire <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u16_u1_105_inst flow-through 
    process(UGT_u16_u1_105_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:UGT_u16_u1_105_inst:flowthrough inputs: " & " num_blk_60 = "& Convert_SLV_To_Hex_String(num_blk_60) & " konst_104_wire_constant = "& Convert_SLV_To_Hex_String(konst_104_wire_constant) & " outputs:" & " UGT_u16_u1_105_wire= "  & Convert_SLV_To_Hex_String(UGT_u16_u1_105_wire));
      --
    end process; 
    -- binary operator UGT_u16_u1_105_inst
    process(num_blk_60) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_60, konst_104_wire_constant, tmp_var);
      UGT_u16_u1_105_wire <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u16_u1_112_inst flow-through 
    process(UGT_u16_u1_112_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:UGT_u16_u1_112_inst:flowthrough inputs: " & " num_blk_60 = "& Convert_SLV_To_Hex_String(num_blk_60) & " konst_111_wire_constant = "& Convert_SLV_To_Hex_String(konst_111_wire_constant) & " outputs:" & " UGT_u16_u1_112_wire= "  & Convert_SLV_To_Hex_String(UGT_u16_u1_112_wire));
      --
    end process; 
    -- binary operator UGT_u16_u1_112_inst
    process(num_blk_60) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_60, konst_111_wire_constant, tmp_var);
      UGT_u16_u1_112_wire <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u16_u1_126_inst flow-through 
    process(c4_127) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:UGT_u16_u1_126_inst:flowthrough inputs: " & " ADD_u16_u16_124_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_124_wire) & " konst_125_wire_constant = "& Convert_SLV_To_Hex_String(konst_125_wire_constant) & " outputs:" & " c4_127= "  & Convert_SLV_To_Hex_String(c4_127));
      --
    end process; 
    -- binary operator UGT_u16_u1_126_inst
    process(ADD_u16_u16_124_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_124_wire, konst_125_wire_constant, tmp_var);
      c4_127 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u16_u1_294_inst flow-through 
    process(UGT_u16_u1_294_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:UGT_u16_u1_294_inst:flowthrough inputs: " & " ADD_u16_u16_292_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_292_wire) & " konst_293_wire_constant = "& Convert_SLV_To_Hex_String(konst_293_wire_constant) & " outputs:" & " UGT_u16_u1_294_wire= "  & Convert_SLV_To_Hex_String(UGT_u16_u1_294_wire));
      --
    end process; 
    -- binary operator UGT_u16_u1_294_inst
    process(ADD_u16_u16_292_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_292_wire, konst_293_wire_constant, tmp_var);
      UGT_u16_u1_294_wire <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u16_u1_92_inst flow-through 
    process(UGT_u16_u1_92_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:UGT_u16_u1_92_inst:flowthrough inputs: " & " num_blk_60 = "& Convert_SLV_To_Hex_String(num_blk_60) & " konst_91_wire_constant = "& Convert_SLV_To_Hex_String(konst_91_wire_constant) & " outputs:" & " UGT_u16_u1_92_wire= "  & Convert_SLV_To_Hex_String(UGT_u16_u1_92_wire));
      --
    end process; 
    -- binary operator UGT_u16_u1_92_inst
    process(num_blk_60) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_60, konst_91_wire_constant, tmp_var);
      UGT_u16_u1_92_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u16_u1_302_inst flow-through 
    process(ULT_u16_u1_302_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ULT_u16_u1_302_inst:flowthrough inputs: " & " n_left_287 = "& Convert_SLV_To_Hex_String(n_left_287) & " konst_301_wire_constant = "& Convert_SLV_To_Hex_String(konst_301_wire_constant) & " outputs:" & " ULT_u16_u1_302_wire= "  & Convert_SLV_To_Hex_String(ULT_u16_u1_302_wire));
      --
    end process; 
    -- binary operator ULT_u16_u1_302_inst
    process(n_left_287) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_left_287, konst_301_wire_constant, tmp_var);
      ULT_u16_u1_302_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u16_u1_38_inst flow-through 
    process(ULT_u16_u1_38_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ULT_u16_u1_38_inst:flowthrough inputs: " & " num_cont_buffer = "& Convert_SLV_To_Hex_String(num_cont_buffer) & " konst_37_wire_constant = "& Convert_SLV_To_Hex_String(konst_37_wire_constant) & " outputs:" & " ULT_u16_u1_38_wire= "  & Convert_SLV_To_Hex_String(ULT_u16_u1_38_wire));
      --
    end process; 
    -- binary operator ULT_u16_u1_38_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(num_cont_buffer, konst_37_wire_constant, tmp_var);
      ULT_u16_u1_38_wire <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_132_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_132_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:array_obj_ref_132_index_offset:started:   inputs: " & " R_address_131_scaled = "& Convert_SLV_To_Hex_String(R_address_131_scaled) & " array_obj_ref_132_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_132_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_132_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:array_obj_ref_132_index_offset:finished:  outputs: " & " array_obj_ref_132_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_132_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (42) : array_obj_ref_132_index_offset 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_131_scaled;
      array_obj_ref_132_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_132_index_offset_req_0;
      array_obj_ref_132_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_132_index_offset_req_1;
      array_obj_ref_132_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- logger for split-operator ptr_deref_137_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_137_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ptr_deref_137_load_0:started:   inputs: " & " ptr_deref_137_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_137_word_address_0));
          --
        end if; 
        if ptr_deref_137_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:ptr_deref_137_load_0:finished:  outputs: " & " ptr_deref_137_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_137_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : ptr_deref_137_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_137_load_0_req_0,
        ptr_deref_137_load_0_ack_0,
        ptr_deref_137_load_0_req_1,
        ptr_deref_137_load_0_ack_1,
        "ptr_deref_137_load_0",
        "memory_space_1" ,
        ptr_deref_137_data_0,
        ptr_deref_137_word_address_0,
        "ptr_deref_137_data_0",
        "ptr_deref_137_word_address_0" -- 
      );
      reqL_unguarded(0) <= ptr_deref_137_load_0_req_0;
      ptr_deref_137_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_137_load_0_req_1;
      ptr_deref_137_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_137_word_address_0;
      ptr_deref_137_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator WPIPE_input_pipe1_166_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_input_pipe1_166_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:WPIPE_input_pipe1_166_inst:started:   PipeWrite to input_pipe1 inputs: " & " c2_159_delayed_14_0_164 (guard)= " & Convert_SLV_To_String(c2_159_delayed_14_0_164) & " w2_146 = "& Convert_SLV_To_Hex_String(w2_146));
          --
        end if; 
        if WPIPE_input_pipe1_166_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:WPIPE_input_pipe1_166_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator WPIPE_input_pipe1_159_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_input_pipe1_159_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:WPIPE_input_pipe1_159_inst:started:   PipeWrite to input_pipe1 inputs: " & " c1_155_delayed_14_0_157 (guard)= " & Convert_SLV_To_String(c1_155_delayed_14_0_157) & " w1_142 = "& Convert_SLV_To_Hex_String(w1_142));
          --
        end if; 
        if WPIPE_input_pipe1_159_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:WPIPE_input_pipe1_159_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator WPIPE_input_pipe1_173_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_input_pipe1_173_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:WPIPE_input_pipe1_173_inst:started:   PipeWrite to input_pipe1 inputs: " & " c3_163_delayed_14_0_171 (guard)= " & Convert_SLV_To_String(c3_163_delayed_14_0_171) & " w3_150 = "& Convert_SLV_To_Hex_String(w3_150));
          --
        end if; 
        if WPIPE_input_pipe1_173_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:WPIPE_input_pipe1_173_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator WPIPE_input_pipe1_180_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_input_pipe1_180_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:WPIPE_input_pipe1_180_inst:started:   PipeWrite to input_pipe1 inputs: " & " c4_167_delayed_14_0_178 (guard)= " & Convert_SLV_To_String(c4_167_delayed_14_0_178) & " w4_154 = "& Convert_SLV_To_Hex_String(w4_154));
          --
        end if; 
        if WPIPE_input_pipe1_180_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:access_T:DP:WPIPE_input_pipe1_180_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_input_pipe1_166_inst WPIPE_input_pipe1_159_inst WPIPE_input_pipe1_173_inst WPIPE_input_pipe1_180_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_input_pipe1_166_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_input_pipe1_159_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_input_pipe1_173_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_input_pipe1_180_inst_req_0;
      WPIPE_input_pipe1_166_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_input_pipe1_159_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_input_pipe1_173_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_input_pipe1_180_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_input_pipe1_166_inst_req_1;
      update_req_unguarded(2) <= WPIPE_input_pipe1_159_inst_req_1;
      update_req_unguarded(1) <= WPIPE_input_pipe1_173_inst_req_1;
      update_req_unguarded(0) <= WPIPE_input_pipe1_180_inst_req_1;
      WPIPE_input_pipe1_166_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_input_pipe1_159_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_input_pipe1_173_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_input_pipe1_180_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= c4_167_delayed_14_0_178(0);
      guard_vector(1)  <= c3_163_delayed_14_0_171(0);
      guard_vector(2)  <= c1_155_delayed_14_0_157(0);
      guard_vector(3)  <= c2_159_delayed_14_0_164(0);
      data_in <= w2_146 & w1_142 & w3_150 & w4_154;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 16, num_reqs => 4, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(95 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(127 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_1120_start: Boolean;
  signal convolution3D_CP_1120_symbol: Boolean;
  -- volatile/operator module components. 
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_529_inst_req_1 : boolean;
  signal type_cast_547_inst_req_0 : boolean;
  signal type_cast_740_inst_ack_0 : boolean;
  signal ptr_deref_652_store_0_req_1 : boolean;
  signal type_cast_470_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_640_inst_req_0 : boolean;
  signal type_cast_608_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_591_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_640_inst_ack_1 : boolean;
  signal type_cast_525_inst_ack_1 : boolean;
  signal if_stmt_666_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_640_inst_req_1 : boolean;
  signal type_cast_525_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_591_inst_ack_1 : boolean;
  signal type_cast_595_inst_ack_1 : boolean;
  signal type_cast_538_inst_ack_1 : boolean;
  signal type_cast_470_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_604_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_591_inst_ack_0 : boolean;
  signal type_cast_529_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_604_inst_req_0 : boolean;
  signal type_cast_470_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_640_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_604_inst_ack_1 : boolean;
  signal type_cast_644_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_604_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_622_inst_ack_1 : boolean;
  signal if_stmt_717_branch_ack_1 : boolean;
  signal addr_of_588_final_reg_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_591_inst_req_1 : boolean;
  signal ptr_deref_652_store_0_req_0 : boolean;
  signal ptr_deref_652_store_0_ack_0 : boolean;
  signal addr_of_588_final_reg_req_0 : boolean;
  signal type_cast_644_inst_req_0 : boolean;
  signal type_cast_547_inst_req_1 : boolean;
  signal addr_of_588_final_reg_ack_0 : boolean;
  signal if_stmt_1055_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_622_inst_ack_0 : boolean;
  signal type_cast_470_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_622_inst_req_0 : boolean;
  signal type_cast_538_inst_req_1 : boolean;
  signal type_cast_525_inst_ack_0 : boolean;
  signal if_stmt_666_branch_req_0 : boolean;
  signal type_cast_595_inst_req_1 : boolean;
  signal if_stmt_666_branch_ack_0 : boolean;
  signal type_cast_552_inst_ack_0 : boolean;
  signal type_cast_547_inst_ack_1 : boolean;
  signal addr_of_588_final_reg_ack_1 : boolean;
  signal type_cast_547_inst_ack_0 : boolean;
  signal type_cast_538_inst_req_0 : boolean;
  signal type_cast_644_inst_req_1 : boolean;
  signal type_cast_595_inst_ack_0 : boolean;
  signal if_stmt_717_branch_ack_0 : boolean;
  signal ptr_deref_652_store_0_ack_1 : boolean;
  signal if_stmt_504_branch_req_0 : boolean;
  signal if_stmt_1106_branch_ack_1 : boolean;
  signal type_cast_538_inst_ack_0 : boolean;
  signal array_obj_ref_587_index_offset_req_0 : boolean;
  signal type_cast_552_inst_req_0 : boolean;
  signal array_obj_ref_587_index_offset_ack_0 : boolean;
  signal type_cast_626_inst_req_0 : boolean;
  signal array_obj_ref_587_index_offset_req_1 : boolean;
  signal array_obj_ref_587_index_offset_ack_1 : boolean;
  signal type_cast_608_inst_req_0 : boolean;
  signal type_cast_626_inst_ack_0 : boolean;
  signal if_stmt_504_branch_ack_1 : boolean;
  signal type_cast_608_inst_ack_0 : boolean;
  signal type_cast_529_inst_ack_0 : boolean;
  signal type_cast_595_inst_req_0 : boolean;
  signal type_cast_740_inst_req_0 : boolean;
  signal type_cast_740_inst_req_1 : boolean;
  signal call_stmt_1232_call_ack_1 : boolean;
  signal type_cast_740_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_760_inst_ack_1 : boolean;
  signal call_stmt_1327_call_ack_1 : boolean;
  signal call_stmt_1360_call_req_1 : boolean;
  signal type_cast_525_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_622_inst_req_1 : boolean;
  signal if_stmt_717_branch_req_0 : boolean;
  signal type_cast_764_inst_ack_0 : boolean;
  signal type_cast_764_inst_req_1 : boolean;
  signal call_stmt_1232_call_req_1 : boolean;
  signal type_cast_764_inst_ack_1 : boolean;
  signal type_cast_1130_inst_req_1 : boolean;
  signal type_cast_1130_inst_ack_1 : boolean;
  signal type_cast_736_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_760_inst_req_0 : boolean;
  signal type_cast_736_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_760_inst_ack_0 : boolean;
  signal type_cast_736_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_760_inst_req_1 : boolean;
  signal call_stmt_1327_call_req_0 : boolean;
  signal phi_stmt_575_ack_0 : boolean;
  signal call_stmt_1327_call_req_1 : boolean;
  signal type_cast_764_inst_req_0 : boolean;
  signal type_cast_736_inst_ack_0 : boolean;
  signal type_cast_529_inst_req_0 : boolean;
  signal type_cast_466_inst_ack_1 : boolean;
  signal addr_of_1222_final_reg_req_0 : boolean;
  signal type_cast_626_inst_ack_1 : boolean;
  signal type_cast_626_inst_req_1 : boolean;
  signal type_cast_552_inst_ack_1 : boolean;
  signal if_stmt_504_branch_ack_0 : boolean;
  signal type_cast_466_inst_req_1 : boolean;
  signal type_cast_552_inst_req_1 : boolean;
  signal type_cast_608_inst_ack_1 : boolean;
  signal type_cast_644_inst_ack_1 : boolean;
  signal if_stmt_1106_branch_ack_0 : boolean;
  signal if_stmt_1055_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1154_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_437_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_437_inst_ack_0 : boolean;
  signal addr_of_1222_final_reg_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_437_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_437_inst_ack_1 : boolean;
  signal type_cast_1364_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_440_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_440_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_440_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_440_inst_ack_1 : boolean;
  signal call_stmt_1327_call_ack_0 : boolean;
  signal call_stmt_1360_call_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_443_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_443_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_443_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_443_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_446_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_446_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_446_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_446_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_449_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_449_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_449_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_449_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_452_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_452_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_452_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_452_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_455_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_455_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_455_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_455_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_458_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_458_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_458_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_458_inst_ack_1 : boolean;
  signal type_cast_462_inst_req_0 : boolean;
  signal type_cast_462_inst_ack_0 : boolean;
  signal type_cast_462_inst_req_1 : boolean;
  signal type_cast_462_inst_ack_1 : boolean;
  signal type_cast_466_inst_req_0 : boolean;
  signal type_cast_466_inst_ack_0 : boolean;
  signal if_stmt_788_branch_req_0 : boolean;
  signal if_stmt_1106_branch_req_0 : boolean;
  signal if_stmt_788_branch_ack_1 : boolean;
  signal if_stmt_788_branch_ack_0 : boolean;
  signal type_cast_1290_inst_ack_1 : boolean;
  signal array_obj_ref_1221_index_offset_ack_1 : boolean;
  signal array_obj_ref_1221_index_offset_req_1 : boolean;
  signal type_cast_1364_inst_ack_0 : boolean;
  signal array_obj_ref_827_index_offset_req_0 : boolean;
  signal array_obj_ref_827_index_offset_ack_0 : boolean;
  signal array_obj_ref_827_index_offset_req_1 : boolean;
  signal call_stmt_1232_call_ack_0 : boolean;
  signal array_obj_ref_827_index_offset_ack_1 : boolean;
  signal call_stmt_1334_call_ack_1 : boolean;
  signal call_stmt_1232_call_req_0 : boolean;
  signal call_stmt_1360_call_ack_0 : boolean;
  signal addr_of_828_final_reg_req_0 : boolean;
  signal addr_of_828_final_reg_ack_0 : boolean;
  signal call_stmt_1360_call_req_0 : boolean;
  signal addr_of_828_final_reg_req_1 : boolean;
  signal addr_of_828_final_reg_ack_1 : boolean;
  signal type_cast_1290_inst_req_1 : boolean;
  signal type_cast_1290_inst_ack_0 : boolean;
  signal type_cast_1290_inst_req_0 : boolean;
  signal ptr_deref_831_store_0_req_0 : boolean;
  signal if_stmt_1182_branch_ack_0 : boolean;
  signal ptr_deref_831_store_0_ack_0 : boolean;
  signal ptr_deref_831_store_0_req_1 : boolean;
  signal ptr_deref_831_store_0_ack_1 : boolean;
  signal type_cast_1323_inst_ack_1 : boolean;
  signal type_cast_1364_inst_req_0 : boolean;
  signal type_cast_838_inst_req_0 : boolean;
  signal type_cast_838_inst_ack_0 : boolean;
  signal type_cast_838_inst_req_1 : boolean;
  signal ptr_deref_1225_store_0_ack_1 : boolean;
  signal type_cast_838_inst_ack_1 : boolean;
  signal phi_stmt_575_req_0 : boolean;
  signal phi_stmt_575_req_1 : boolean;
  signal type_cast_1281_inst_ack_1 : boolean;
  signal if_stmt_1182_branch_ack_1 : boolean;
  signal type_cast_842_inst_req_0 : boolean;
  signal ptr_deref_1225_store_0_req_1 : boolean;
  signal type_cast_842_inst_ack_0 : boolean;
  signal type_cast_842_inst_req_1 : boolean;
  signal type_cast_842_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1371_inst_ack_1 : boolean;
  signal type_cast_581_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1371_inst_req_1 : boolean;
  signal type_cast_1281_inst_req_1 : boolean;
  signal type_cast_846_inst_req_0 : boolean;
  signal type_cast_846_inst_ack_0 : boolean;
  signal type_cast_846_inst_req_1 : boolean;
  signal type_cast_846_inst_ack_1 : boolean;
  signal type_cast_581_inst_req_1 : boolean;
  signal type_cast_1323_inst_req_1 : boolean;
  signal type_cast_1356_inst_ack_1 : boolean;
  signal array_obj_ref_1221_index_offset_ack_0 : boolean;
  signal type_cast_1356_inst_req_1 : boolean;
  signal if_stmt_884_branch_req_0 : boolean;
  signal array_obj_ref_1221_index_offset_req_0 : boolean;
  signal if_stmt_884_branch_ack_1 : boolean;
  signal if_stmt_884_branch_ack_0 : boolean;
  signal type_cast_1281_inst_ack_0 : boolean;
  signal call_stmt_1334_call_req_1 : boolean;
  signal type_cast_1134_inst_ack_1 : boolean;
  signal type_cast_1281_inst_req_0 : boolean;
  signal type_cast_905_inst_req_0 : boolean;
  signal type_cast_905_inst_ack_0 : boolean;
  signal type_cast_1356_inst_ack_0 : boolean;
  signal type_cast_905_inst_req_1 : boolean;
  signal type_cast_905_inst_ack_1 : boolean;
  signal if_stmt_1182_branch_req_0 : boolean;
  signal type_cast_1356_inst_req_0 : boolean;
  signal type_cast_909_inst_req_0 : boolean;
  signal type_cast_909_inst_ack_0 : boolean;
  signal type_cast_909_inst_req_1 : boolean;
  signal ptr_deref_1225_store_0_ack_0 : boolean;
  signal type_cast_909_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1371_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1371_inst_req_0 : boolean;
  signal type_cast_918_inst_req_0 : boolean;
  signal ptr_deref_1225_store_0_req_0 : boolean;
  signal type_cast_918_inst_ack_0 : boolean;
  signal type_cast_1134_inst_req_1 : boolean;
  signal type_cast_918_inst_req_1 : boolean;
  signal type_cast_918_inst_ack_1 : boolean;
  signal type_cast_581_inst_ack_0 : boolean;
  signal type_cast_1271_inst_ack_1 : boolean;
  signal type_cast_1271_inst_req_1 : boolean;
  signal type_cast_927_inst_req_0 : boolean;
  signal type_cast_927_inst_ack_0 : boolean;
  signal type_cast_927_inst_req_1 : boolean;
  signal type_cast_927_inst_ack_1 : boolean;
  signal type_cast_581_inst_req_0 : boolean;
  signal type_cast_1271_inst_ack_0 : boolean;
  signal type_cast_1271_inst_req_0 : boolean;
  signal type_cast_936_inst_req_0 : boolean;
  signal type_cast_936_inst_ack_0 : boolean;
  signal type_cast_936_inst_req_1 : boolean;
  signal type_cast_936_inst_ack_1 : boolean;
  signal if_stmt_1346_branch_ack_0 : boolean;
  signal type_cast_941_inst_req_0 : boolean;
  signal type_cast_941_inst_ack_0 : boolean;
  signal type_cast_941_inst_req_1 : boolean;
  signal type_cast_941_inst_ack_1 : boolean;
  signal type_cast_1323_inst_ack_0 : boolean;
  signal call_stmt_1334_call_ack_0 : boolean;
  signal type_cast_1158_inst_ack_1 : boolean;
  signal type_cast_1158_inst_req_1 : boolean;
  signal type_cast_1323_inst_req_0 : boolean;
  signal array_obj_ref_976_index_offset_req_0 : boolean;
  signal array_obj_ref_976_index_offset_ack_0 : boolean;
  signal type_cast_1130_inst_ack_0 : boolean;
  signal array_obj_ref_976_index_offset_req_1 : boolean;
  signal array_obj_ref_976_index_offset_ack_1 : boolean;
  signal call_stmt_1334_call_req_0 : boolean;
  signal type_cast_1130_inst_req_0 : boolean;
  signal addr_of_977_final_reg_req_0 : boolean;
  signal addr_of_977_final_reg_ack_0 : boolean;
  signal if_stmt_1346_branch_ack_1 : boolean;
  signal addr_of_977_final_reg_req_1 : boolean;
  signal addr_of_977_final_reg_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1247_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_980_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_980_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_980_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_980_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1247_inst_req_1 : boolean;
  signal type_cast_1158_inst_ack_0 : boolean;
  signal type_cast_1158_inst_req_0 : boolean;
  signal type_cast_984_inst_req_0 : boolean;
  signal type_cast_984_inst_ack_0 : boolean;
  signal if_stmt_1055_branch_ack_0 : boolean;
  signal type_cast_984_inst_req_1 : boolean;
  signal type_cast_984_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_993_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_993_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_993_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_993_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1247_inst_ack_0 : boolean;
  signal type_cast_997_inst_req_0 : boolean;
  signal type_cast_997_inst_ack_0 : boolean;
  signal if_stmt_1346_branch_req_0 : boolean;
  signal type_cast_997_inst_req_1 : boolean;
  signal type_cast_997_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1247_inst_req_0 : boolean;
  signal type_cast_1319_inst_ack_1 : boolean;
  signal type_cast_1319_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1011_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1011_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1011_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1011_inst_ack_1 : boolean;
  signal type_cast_1015_inst_req_0 : boolean;
  signal type_cast_1015_inst_ack_0 : boolean;
  signal type_cast_1015_inst_req_1 : boolean;
  signal type_cast_1015_inst_ack_1 : boolean;
  signal type_cast_1319_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1029_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1029_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1029_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1029_inst_ack_1 : boolean;
  signal type_cast_1033_inst_req_0 : boolean;
  signal type_cast_1033_inst_ack_0 : boolean;
  signal type_cast_1033_inst_req_1 : boolean;
  signal type_cast_1033_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1244_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1244_inst_req_1 : boolean;
  signal WPIPE_num_out_pipe_1244_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_1244_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1154_inst_ack_1 : boolean;
  signal addr_of_1222_final_reg_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1154_inst_req_1 : boolean;
  signal addr_of_1222_final_reg_req_1 : boolean;
  signal type_cast_1319_inst_req_0 : boolean;
  signal type_cast_1134_inst_ack_0 : boolean;
  signal ptr_deref_1041_store_0_req_0 : boolean;
  signal ptr_deref_1041_store_0_ack_0 : boolean;
  signal type_cast_1134_inst_req_0 : boolean;
  signal ptr_deref_1041_store_0_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1154_inst_ack_0 : boolean;
  signal ptr_deref_1041_store_0_ack_1 : boolean;
  signal type_cast_1364_inst_ack_1 : boolean;
  signal phi_stmt_697_req_1 : boolean;
  signal type_cast_700_inst_req_0 : boolean;
  signal type_cast_700_inst_ack_0 : boolean;
  signal type_cast_700_inst_req_1 : boolean;
  signal type_cast_700_inst_ack_1 : boolean;
  signal phi_stmt_697_req_0 : boolean;
  signal phi_stmt_697_ack_0 : boolean;
  signal type_cast_747_inst_req_0 : boolean;
  signal type_cast_747_inst_ack_0 : boolean;
  signal type_cast_747_inst_req_1 : boolean;
  signal type_cast_747_inst_ack_1 : boolean;
  signal phi_stmt_744_req_0 : boolean;
  signal type_cast_754_inst_req_0 : boolean;
  signal type_cast_754_inst_ack_0 : boolean;
  signal type_cast_754_inst_req_1 : boolean;
  signal type_cast_754_inst_ack_1 : boolean;
  signal phi_stmt_751_req_0 : boolean;
  signal phi_stmt_744_req_1 : boolean;
  signal phi_stmt_751_req_1 : boolean;
  signal phi_stmt_744_ack_0 : boolean;
  signal phi_stmt_751_ack_0 : boolean;
  signal type_cast_798_inst_req_0 : boolean;
  signal type_cast_798_inst_ack_0 : boolean;
  signal type_cast_798_inst_req_1 : boolean;
  signal type_cast_798_inst_ack_1 : boolean;
  signal phi_stmt_795_req_0 : boolean;
  signal phi_stmt_795_ack_0 : boolean;
  signal phi_stmt_964_req_0 : boolean;
  signal type_cast_970_inst_req_0 : boolean;
  signal type_cast_970_inst_ack_0 : boolean;
  signal type_cast_970_inst_req_1 : boolean;
  signal type_cast_970_inst_ack_1 : boolean;
  signal phi_stmt_964_req_1 : boolean;
  signal phi_stmt_964_ack_0 : boolean;
  signal type_cast_1089_inst_req_0 : boolean;
  signal type_cast_1089_inst_ack_0 : boolean;
  signal type_cast_1089_inst_req_1 : boolean;
  signal type_cast_1089_inst_ack_1 : boolean;
  signal phi_stmt_1086_req_0 : boolean;
  signal phi_stmt_1086_req_1 : boolean;
  signal phi_stmt_1086_ack_0 : boolean;
  signal type_cast_1141_inst_req_0 : boolean;
  signal type_cast_1141_inst_ack_0 : boolean;
  signal type_cast_1141_inst_req_1 : boolean;
  signal type_cast_1141_inst_ack_1 : boolean;
  signal phi_stmt_1138_req_0 : boolean;
  signal type_cast_1148_inst_req_0 : boolean;
  signal type_cast_1148_inst_ack_0 : boolean;
  signal type_cast_1148_inst_req_1 : boolean;
  signal type_cast_1148_inst_ack_1 : boolean;
  signal phi_stmt_1145_req_0 : boolean;
  signal phi_stmt_1138_req_1 : boolean;
  signal phi_stmt_1145_req_1 : boolean;
  signal phi_stmt_1138_ack_0 : boolean;
  signal phi_stmt_1145_ack_0 : boolean;
  signal type_cast_1192_inst_req_0 : boolean;
  signal type_cast_1192_inst_ack_0 : boolean;
  signal type_cast_1192_inst_req_1 : boolean;
  signal type_cast_1192_inst_ack_1 : boolean;
  signal phi_stmt_1189_req_0 : boolean;
  signal phi_stmt_1189_ack_0 : boolean;
  signal phi_stmt_1299_req_1 : boolean;
  signal type_cast_1302_inst_req_0 : boolean;
  signal type_cast_1302_inst_ack_0 : boolean;
  signal type_cast_1302_inst_req_1 : boolean;
  signal type_cast_1302_inst_ack_1 : boolean;
  signal phi_stmt_1299_req_0 : boolean;
  signal phi_stmt_1299_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_1120_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1120_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_1120_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1120_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,convolution3D_CP_1120_start,"convolution3D cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,convolution3D_CP_1120_symbol, "convolution3D cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_1120: Block -- control-path 
    signal convolution3D_CP_1120_elements: BooleanArray(249 downto 0);
    -- 
  begin -- 
    convolution3D_CP_1120_elements(0) <= convolution3D_CP_1120_start;
    convolution3D_CP_1120_symbol <= convolution3D_CP_1120_elements(181);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	18 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	22 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_470_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_470_update_start_
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_470_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_466_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_435/$entry
      -- CP-element group 0: 	 branch_block_stmt_435/branch_block_stmt_435__entry__
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503__entry__
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/$entry
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_437_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_437_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_437_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_462_update_start_
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_462_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_462_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_466_update_start_
      -- CP-element group 0: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_466_Update/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_470_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_466_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_437_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_462_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_470_inst_req_1); -- 
    cr_1367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_466_inst_req_1); -- 
    rr_1236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => RPIPE_maxpool_input_pipe_437_inst_req_0); -- 
    cr_1353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_462_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_437_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_437_update_start_
      -- CP-element group 1: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_437_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_437_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_437_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_437_Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_437_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_437_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_1237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_437_inst_ack_0, ack => convolution3D_CP_1120_elements(1)); -- 
    cr_1241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(1), ack => RPIPE_maxpool_input_pipe_437_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	17 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_437_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_437_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_437_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_440_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_440_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_440_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_462_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_462_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_462_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_437_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_440_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_462_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_437_inst_ack_1, ack => convolution3D_CP_1120_elements(2)); -- 
    rr_1250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(2), ack => RPIPE_maxpool_input_pipe_440_inst_req_0); -- 
    rr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(2), ack => type_cast_462_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_440_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_440_update_start_
      -- CP-element group 3: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_440_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_440_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_440_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_440_Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_440_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_440_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_1251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_440_inst_ack_0, ack => convolution3D_CP_1120_elements(3)); -- 
    cr_1255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(3), ack => RPIPE_maxpool_input_pipe_440_inst_req_1); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	19 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_440_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_440_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_440_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_443_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_443_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_443_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_466_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_466_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_466_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_440_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_443_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_466_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_440_inst_ack_1, ack => convolution3D_CP_1120_elements(4)); -- 
    rr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(4), ack => RPIPE_maxpool_input_pipe_443_inst_req_0); -- 
    rr_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(4), ack => type_cast_466_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_443_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_443_update_start_
      -- CP-element group 5: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_443_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_443_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_443_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_443_Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_443_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_443_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_443_inst_ack_0, ack => convolution3D_CP_1120_elements(5)); -- 
    cr_1269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(5), ack => RPIPE_maxpool_input_pipe_443_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	21 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_470_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_470_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_470_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_443_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_443_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_443_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_446_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_446_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_446_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_443_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_446_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_470_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_443_inst_ack_1, ack => convolution3D_CP_1120_elements(6)); -- 
    rr_1278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(6), ack => RPIPE_maxpool_input_pipe_446_inst_req_0); -- 
    rr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(6), ack => type_cast_470_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_446_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_446_update_start_
      -- CP-element group 7: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_446_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_446_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_446_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_446_Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_446_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_446_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_1279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_446_inst_ack_0, ack => convolution3D_CP_1120_elements(7)); -- 
    cr_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(7), ack => RPIPE_maxpool_input_pipe_446_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_446_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_446_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_446_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_449_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_449_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_449_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_446_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_449_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_446_inst_ack_1, ack => convolution3D_CP_1120_elements(8)); -- 
    rr_1292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(8), ack => RPIPE_maxpool_input_pipe_449_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_449_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_449_update_start_
      -- CP-element group 9: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_449_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_449_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_449_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_449_Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_449_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_449_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_449_inst_ack_0, ack => convolution3D_CP_1120_elements(9)); -- 
    cr_1297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(9), ack => RPIPE_maxpool_input_pipe_449_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_449_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_449_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_449_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_452_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_452_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_452_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_449_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_452_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_449_inst_ack_1, ack => convolution3D_CP_1120_elements(10)); -- 
    rr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(10), ack => RPIPE_maxpool_input_pipe_452_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_452_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_452_update_start_
      -- CP-element group 11: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_452_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_452_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_452_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_452_Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_452_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_452_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_452_inst_ack_0, ack => convolution3D_CP_1120_elements(11)); -- 
    cr_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(11), ack => RPIPE_maxpool_input_pipe_452_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_452_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_452_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_452_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_455_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_455_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_455_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_452_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_455_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_452_inst_ack_1, ack => convolution3D_CP_1120_elements(12)); -- 
    rr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(12), ack => RPIPE_maxpool_input_pipe_455_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_455_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_455_update_start_
      -- CP-element group 13: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_455_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_455_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_455_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_455_Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_455_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_455_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_455_inst_ack_0, ack => convolution3D_CP_1120_elements(13)); -- 
    cr_1325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(13), ack => RPIPE_maxpool_input_pipe_455_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_455_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_455_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_455_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_458_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_458_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_458_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_455_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_458_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_455_inst_ack_1, ack => convolution3D_CP_1120_elements(14)); -- 
    rr_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(14), ack => RPIPE_maxpool_input_pipe_458_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_458_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_458_update_start_
      -- CP-element group 15: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_458_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_458_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_458_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_458_Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_458_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_458_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_458_inst_ack_0, ack => convolution3D_CP_1120_elements(15)); -- 
    cr_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(15), ack => RPIPE_maxpool_input_pipe_458_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	23 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_458_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_458_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/RPIPE_maxpool_input_pipe_458_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_458_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_458_inst_ack_1, ack => convolution3D_CP_1120_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_462_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_462_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_462_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_462_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_462_inst_ack_0, ack => convolution3D_CP_1120_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	0 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	23 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_462_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_462_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_462_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_462_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_462_inst_ack_1, ack => convolution3D_CP_1120_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	4 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_466_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_466_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_466_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_466_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_466_inst_ack_0, ack => convolution3D_CP_1120_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	23 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_466_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_466_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_466_Update/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_466_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_466_inst_ack_1, ack => convolution3D_CP_1120_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	6 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_470_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_470_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_470_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_470_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_470_inst_ack_0, ack => convolution3D_CP_1120_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	0 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_470_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_470_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/type_cast_470_Update/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_470_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_470_inst_ack_1, ack => convolution3D_CP_1120_elements(22)); -- 
    -- CP-element group 23:  branch  join  transition  place  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	16 
    -- CP-element group 23: 	18 
    -- CP-element group 23: 	20 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (10) 
      -- CP-element group 23: 	 branch_block_stmt_435/if_stmt_504_eval_test/$entry
      -- CP-element group 23: 	 branch_block_stmt_435/if_stmt_504_if_link/$entry
      -- CP-element group 23: 	 branch_block_stmt_435/if_stmt_504_dead_link/$entry
      -- CP-element group 23: 	 branch_block_stmt_435/if_stmt_504_eval_test/$exit
      -- CP-element group 23: 	 branch_block_stmt_435/if_stmt_504_eval_test/branch_req
      -- CP-element group 23: 	 branch_block_stmt_435/if_stmt_504_else_link/$entry
      -- CP-element group 23: 	 branch_block_stmt_435/R_cmp195_505_place
      -- CP-element group 23: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503__exit__
      -- CP-element group 23: 	 branch_block_stmt_435/if_stmt_504__entry__
      -- CP-element group 23: 	 branch_block_stmt_435/assign_stmt_438_to_assign_stmt_503/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_504_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(23), ack => if_stmt_504_branch_req_0); -- 
    convolution3D_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(16) & convolution3D_CP_1120_elements(18) & convolution3D_CP_1120_elements(20) & convolution3D_CP_1120_elements(22);
      gj_convolution3D_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	29 
    -- CP-element group 24: 	30 
    -- CP-element group 24: 	31 
    -- CP-element group 24: 	34 
    -- CP-element group 24: 	36 
    -- CP-element group 24:  members (36) 
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_529_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_525_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_529_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_529_update_start_
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_552_update_start_
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_547_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_538_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_538_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_538_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_538_update_start_
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_547_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_525_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_529_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_538_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_538_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_435/if_stmt_504_if_link/$exit
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_547_update_start_
      -- CP-element group 24: 	 branch_block_stmt_435/if_stmt_504_if_link/if_choice_transition
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_525_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_435/entry_bbx_xnph197_PhiReq/$entry
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_525_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_525_update_start_
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_525_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_529_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_435/merge_stmt_510_PhiAck/dummy
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/$entry
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_529_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_435/entry_bbx_xnph197
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_552_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_552_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_435/merge_stmt_510__exit__
      -- CP-element group 24: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572__entry__
      -- CP-element group 24: 	 branch_block_stmt_435/merge_stmt_510_PhiAck/$exit
      -- CP-element group 24: 	 branch_block_stmt_435/merge_stmt_510_PhiAck/$entry
      -- CP-element group 24: 	 branch_block_stmt_435/merge_stmt_510_PhiReqMerge
      -- CP-element group 24: 	 branch_block_stmt_435/entry_bbx_xnph197_PhiReq/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_504_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_529_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_525_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_547_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_538_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_538_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_525_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_529_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_552_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_1395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_504_branch_ack_1, ack => convolution3D_CP_1120_elements(24)); -- 
    cr_1431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(24), ack => type_cast_529_inst_req_1); -- 
    cr_1417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(24), ack => type_cast_525_inst_req_1); -- 
    cr_1459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(24), ack => type_cast_547_inst_req_1); -- 
    cr_1445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(24), ack => type_cast_538_inst_req_1); -- 
    rr_1440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(24), ack => type_cast_538_inst_req_0); -- 
    rr_1412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(24), ack => type_cast_525_inst_req_0); -- 
    rr_1426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(24), ack => type_cast_529_inst_req_0); -- 
    cr_1473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(24), ack => type_cast_552_inst_req_1); -- 
    -- CP-element group 25:  transition  place  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	188 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_435/if_stmt_504_else_link/$exit
      -- CP-element group 25: 	 branch_block_stmt_435/entry_forx_xend
      -- CP-element group 25: 	 branch_block_stmt_435/if_stmt_504_else_link/else_choice_transition
      -- CP-element group 25: 	 branch_block_stmt_435/entry_forx_xend_PhiReq/$entry
      -- CP-element group 25: 	 branch_block_stmt_435/entry_forx_xend_PhiReq/phi_stmt_697/$entry
      -- CP-element group 25: 	 branch_block_stmt_435/entry_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_504_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_1399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_504_branch_ack_0, ack => convolution3D_CP_1120_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_525_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_525_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_525_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_525_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_525_inst_ack_0, ack => convolution3D_CP_1120_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	32 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_525_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_525_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_525_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_525_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_525_inst_ack_1, ack => convolution3D_CP_1120_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_529_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_529_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_529_Sample/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_529_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_529_inst_ack_0, ack => convolution3D_CP_1120_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_529_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_529_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_529_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_529_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_529_inst_ack_1, ack => convolution3D_CP_1120_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_538_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_538_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_538_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_538_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_0, ack => convolution3D_CP_1120_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	24 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_538_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_538_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_538_Update/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_538_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_1, ack => convolution3D_CP_1120_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	27 
    -- CP-element group 32: 	29 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_547_Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_547_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_547_Sample/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_547_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(32), ack => type_cast_547_inst_req_0); -- 
    convolution3D_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(27) & convolution3D_CP_1120_elements(29) & convolution3D_CP_1120_elements(31);
      gj_convolution3D_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_547_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_547_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_547_Sample/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_547_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_547_inst_ack_0, ack => convolution3D_CP_1120_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	24 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_552_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_552_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_547_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_547_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_552_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_547_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_547_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_552_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_547_inst_ack_1, ack => convolution3D_CP_1120_elements(34)); -- 
    rr_1468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(34), ack => type_cast_552_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_552_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_552_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_552_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_552_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_552_inst_ack_0, ack => convolution3D_CP_1120_elements(35)); -- 
    -- CP-element group 36:  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	24 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	182 
    -- CP-element group 36:  members (9) 
      -- CP-element group 36: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_552_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/$exit
      -- CP-element group 36: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_552_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572/type_cast_552_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_435/assign_stmt_516_to_assign_stmt_572__exit__
      -- CP-element group 36: 	 branch_block_stmt_435/bbx_xnph197_forx_xbody
      -- CP-element group 36: 	 branch_block_stmt_435/bbx_xnph197_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/$entry
      -- CP-element group 36: 	 branch_block_stmt_435/bbx_xnph197_forx_xbody_PhiReq/phi_stmt_575/$entry
      -- CP-element group 36: 	 branch_block_stmt_435/bbx_xnph197_forx_xbody_PhiReq/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_552_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_552_inst_ack_1, ack => convolution3D_CP_1120_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	187 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	60 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_final_index_sum_regn_sample_complete
      -- CP-element group 37: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_final_index_sum_regn_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_587_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_587_index_offset_ack_0, ack => convolution3D_CP_1120_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	187 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (11) 
      -- CP-element group 38: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_offset_calculated
      -- CP-element group 38: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_root_address_calculated
      -- CP-element group 38: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/addr_of_588_request/req
      -- CP-element group 38: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/addr_of_588_request/$entry
      -- CP-element group 38: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_final_index_sum_regn_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_final_index_sum_regn_Update/ack
      -- CP-element group 38: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_base_plus_offset/$entry
      -- CP-element group 38: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_base_plus_offset/sum_rename_ack
      -- CP-element group 38: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/addr_of_588_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_base_plus_offset/sum_rename_req
      -- CP-element group 38: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_base_plus_offset/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_587_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_588_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_587_index_offset_ack_1, ack => convolution3D_CP_1120_elements(38)); -- 
    req_1517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(38), ack => addr_of_588_final_reg_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/addr_of_588_request/$exit
      -- CP-element group 39: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/addr_of_588_request/ack
      -- CP-element group 39: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/addr_of_588_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_588_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_588_final_reg_ack_0, ack => convolution3D_CP_1120_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	187 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	57 
    -- CP-element group 40:  members (19) 
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_word_addrgen/$exit
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_word_addrgen/$entry
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_base_addr_resize/base_resize_ack
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_base_plus_offset/$entry
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_base_addr_resize/$exit
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_base_addr_resize/base_resize_req
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_base_plus_offset/sum_rename_req
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_base_plus_offset/sum_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_base_plus_offset/$exit
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/addr_of_588_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/addr_of_588_complete/$exit
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/addr_of_588_complete/ack
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_base_addr_resize/$entry
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_base_address_resized
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_word_addrgen/root_register_req
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_word_addrgen/root_register_ack
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_root_address_calculated
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_word_address_calculated
      -- CP-element group 40: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_base_address_calculated
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_588_final_reg_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_588_final_reg_ack_1, ack => convolution3D_CP_1120_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	187 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_591_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_591_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_591_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_591_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_591_update_start_
      -- CP-element group 41: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_591_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_591_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_591_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_1532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_591_inst_ack_0, ack => convolution3D_CP_1120_elements(41)); -- 
    cr_1536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(41), ack => RPIPE_maxpool_input_pipe_591_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_591_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_604_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_604_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_591_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_595_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_604_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_595_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_595_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_591_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_591_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_595_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_604_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_591_inst_ack_1, ack => convolution3D_CP_1120_elements(42)); -- 
    rr_1545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(42), ack => type_cast_595_inst_req_0); -- 
    rr_1559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(42), ack => RPIPE_maxpool_input_pipe_604_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_595_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_595_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_595_Sample/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_595_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_595_inst_ack_0, ack => convolution3D_CP_1120_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	187 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	57 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_595_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_595_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_595_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_595_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_595_inst_ack_1, ack => convolution3D_CP_1120_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_604_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_604_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_604_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_604_Update/cr
      -- CP-element group 45: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_604_update_start_
      -- CP-element group 45: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_604_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_604_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_604_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_1560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_604_inst_ack_0, ack => convolution3D_CP_1120_elements(45)); -- 
    cr_1564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(45), ack => RPIPE_maxpool_input_pipe_604_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_604_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_608_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_604_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_604_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_622_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_608_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_608_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_622_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_622_sample_start_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_604_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_608_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_622_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_604_inst_ack_1, ack => convolution3D_CP_1120_elements(46)); -- 
    rr_1573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(46), ack => type_cast_608_inst_req_0); -- 
    rr_1587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(46), ack => RPIPE_maxpool_input_pipe_622_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_608_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_608_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_608_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_608_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_0, ack => convolution3D_CP_1120_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	187 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	57 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_608_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_608_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_608_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_608_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_1, ack => convolution3D_CP_1120_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_622_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_622_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_622_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_622_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_622_update_start_
      -- CP-element group 49: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_622_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_622_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_622_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_1588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_622_inst_ack_0, ack => convolution3D_CP_1120_elements(49)); -- 
    cr_1592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(49), ack => RPIPE_maxpool_input_pipe_622_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_640_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_640_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_622_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_626_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_622_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_626_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_626_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_622_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_640_sample_start_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_622_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_626_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_640_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_622_inst_ack_1, ack => convolution3D_CP_1120_elements(50)); -- 
    rr_1601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(50), ack => type_cast_626_inst_req_0); -- 
    rr_1615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(50), ack => RPIPE_maxpool_input_pipe_640_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_626_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_626_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_626_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_626_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_626_inst_ack_0, ack => convolution3D_CP_1120_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	187 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	57 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_626_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_626_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_626_Update/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_626_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_626_inst_ack_1, ack => convolution3D_CP_1120_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_640_Update/cr
      -- CP-element group 53: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_640_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_640_update_start_
      -- CP-element group 53: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_640_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_640_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_640_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_640_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_640_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_1616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_640_inst_ack_0, ack => convolution3D_CP_1120_elements(53)); -- 
    cr_1620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(53), ack => RPIPE_maxpool_input_pipe_640_inst_req_1); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_640_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_644_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_640_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_644_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_640_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_644_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_640_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_644_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_640_inst_ack_1, ack => convolution3D_CP_1120_elements(54)); -- 
    rr_1629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(54), ack => type_cast_644_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_644_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_644_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_644_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_644_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_644_inst_ack_0, ack => convolution3D_CP_1120_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	187 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_644_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_644_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_644_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_644_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_644_inst_ack_1, ack => convolution3D_CP_1120_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	40 
    -- CP-element group 57: 	44 
    -- CP-element group 57: 	48 
    -- CP-element group 57: 	52 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Sample/word_access_start/$entry
      -- CP-element group 57: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Sample/ptr_deref_652_Split/split_ack
      -- CP-element group 57: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Sample/word_access_start/word_0/rr
      -- CP-element group 57: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Sample/word_access_start/word_0/$entry
      -- CP-element group 57: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Sample/ptr_deref_652_Split/split_req
      -- CP-element group 57: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Sample/ptr_deref_652_Split/$exit
      -- CP-element group 57: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Sample/ptr_deref_652_Split/$entry
      -- CP-element group 57: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_sample_start_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_652_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(57), ack => ptr_deref_652_store_0_req_0); -- 
    convolution3D_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(40) & convolution3D_CP_1120_elements(44) & convolution3D_CP_1120_elements(48) & convolution3D_CP_1120_elements(52) & convolution3D_CP_1120_elements(56);
      gj_convolution3D_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (5) 
      -- CP-element group 58: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Sample/word_access_start/$exit
      -- CP-element group 58: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Sample/word_access_start/word_0/ra
      -- CP-element group 58: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Sample/word_access_start/word_0/$exit
      -- CP-element group 58: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Sample/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_652_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_652_store_0_ack_0, ack => convolution3D_CP_1120_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	187 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Update/word_access_complete/word_0/$exit
      -- CP-element group 59: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Update/word_access_complete/$exit
      -- CP-element group 59: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Update/word_access_complete/word_0/ca
      -- CP-element group 59: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_652_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_652_store_0_ack_1, ack => convolution3D_CP_1120_elements(59)); -- 
    -- CP-element group 60:  branch  join  transition  place  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	37 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (10) 
      -- CP-element group 60: 	 branch_block_stmt_435/if_stmt_666_else_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_435/if_stmt_666_eval_test/$exit
      -- CP-element group 60: 	 branch_block_stmt_435/if_stmt_666_eval_test/$entry
      -- CP-element group 60: 	 branch_block_stmt_435/if_stmt_666_if_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_435/R_exitcond37_667_place
      -- CP-element group 60: 	 branch_block_stmt_435/if_stmt_666_eval_test/branch_req
      -- CP-element group 60: 	 branch_block_stmt_435/if_stmt_666_dead_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/$exit
      -- CP-element group 60: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665__exit__
      -- CP-element group 60: 	 branch_block_stmt_435/if_stmt_666__entry__
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_666_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(60), ack => if_stmt_666_branch_req_0); -- 
    convolution3D_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(37) & convolution3D_CP_1120_elements(59);
      gj_convolution3D_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	189 
    -- CP-element group 61: 	190 
    -- CP-element group 61:  members (24) 
      -- CP-element group 61: 	 branch_block_stmt_435/if_stmt_666_if_link/if_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_435/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 61: 	 branch_block_stmt_435/if_stmt_666_if_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_435/assign_stmt_679_to_assign_stmt_694/$entry
      -- CP-element group 61: 	 branch_block_stmt_435/assign_stmt_679_to_assign_stmt_694/$exit
      -- CP-element group 61: 	 branch_block_stmt_435/merge_stmt_672__exit__
      -- CP-element group 61: 	 branch_block_stmt_435/assign_stmt_679_to_assign_stmt_694__entry__
      -- CP-element group 61: 	 branch_block_stmt_435/assign_stmt_679_to_assign_stmt_694__exit__
      -- CP-element group 61: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 61: 	 branch_block_stmt_435/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_435/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 61: 	 branch_block_stmt_435/merge_stmt_672_PhiReqMerge
      -- CP-element group 61: 	 branch_block_stmt_435/merge_stmt_672_PhiAck/$entry
      -- CP-element group 61: 	 branch_block_stmt_435/merge_stmt_672_PhiAck/$exit
      -- CP-element group 61: 	 branch_block_stmt_435/merge_stmt_672_PhiAck/dummy
      -- CP-element group 61: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/$entry
      -- CP-element group 61: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/type_cast_700/$entry
      -- CP-element group 61: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/type_cast_700/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/type_cast_700/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/type_cast_700/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/type_cast_700/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/type_cast_700/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_666_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_700_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_700_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_666_branch_ack_1, ack => convolution3D_CP_1120_elements(61)); -- 
    rr_2821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(61), ack => type_cast_700_inst_req_0); -- 
    cr_2826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(61), ack => type_cast_700_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	183 
    -- CP-element group 62: 	184 
    -- CP-element group 62:  members (12) 
      -- CP-element group 62: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/type_cast_581/$entry
      -- CP-element group 62: 	 branch_block_stmt_435/if_stmt_666_else_link/$exit
      -- CP-element group 62: 	 branch_block_stmt_435/if_stmt_666_else_link/else_choice_transition
      -- CP-element group 62: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/$entry
      -- CP-element group 62: 	 branch_block_stmt_435/forx_xbody_forx_xbody
      -- CP-element group 62: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/type_cast_581/SplitProtocol/Update/cr
      -- CP-element group 62: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/$entry
      -- CP-element group 62: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/type_cast_581/SplitProtocol/Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/type_cast_581/SplitProtocol/Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/type_cast_581/SplitProtocol/Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 62: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/type_cast_581/SplitProtocol/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_666_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_581_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_581_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_1702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_666_branch_ack_0, ack => convolution3D_CP_1120_elements(62)); -- 
    cr_2772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(62), ack => type_cast_581_inst_req_1); -- 
    rr_2767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(62), ack => type_cast_581_inst_req_0); -- 
    -- CP-element group 63:  transition  place  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	193 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	212 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_435/if_stmt_717_if_link/if_choice_transition
      -- CP-element group 63: 	 branch_block_stmt_435/if_stmt_717_if_link/$exit
      -- CP-element group 63: 	 branch_block_stmt_435/forx_xend_ifx_xend
      -- CP-element group 63: 	 branch_block_stmt_435/forx_xend_ifx_xend_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_435/forx_xend_ifx_xend_PhiReq/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_717_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_1723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_717_branch_ack_1, ack => convolution3D_CP_1120_elements(63)); -- 
    -- CP-element group 64:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	193 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	66 
    -- CP-element group 64: 	68 
    -- CP-element group 64:  members (21) 
      -- CP-element group 64: 	 branch_block_stmt_435/if_stmt_717_else_link/else_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_740_Update/cr
      -- CP-element group 64: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/$entry
      -- CP-element group 64: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_740_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_435/if_stmt_717_else_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_736_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_736_Update/cr
      -- CP-element group 64: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_740_update_start_
      -- CP-element group 64: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_736_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_736_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_736_update_start_
      -- CP-element group 64: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_736_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_435/forx_xend_forx_xbodyx_xix_xpreheader
      -- CP-element group 64: 	 branch_block_stmt_435/merge_stmt_723__exit__
      -- CP-element group 64: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741__entry__
      -- CP-element group 64: 	 branch_block_stmt_435/forx_xend_forx_xbodyx_xix_xpreheader_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_435/forx_xend_forx_xbodyx_xix_xpreheader_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_435/merge_stmt_723_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_435/merge_stmt_723_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_435/merge_stmt_723_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_435/merge_stmt_723_PhiAck/dummy
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_717_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_740_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_736_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_736_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_1727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_717_branch_ack_0, ack => convolution3D_CP_1120_elements(64)); -- 
    cr_1759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(64), ack => type_cast_740_inst_req_1); -- 
    cr_1745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(64), ack => type_cast_736_inst_req_1); -- 
    rr_1740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(64), ack => type_cast_736_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_736_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_736_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_736_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_736_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_736_inst_ack_0, ack => convolution3D_CP_1120_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_740_Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_740_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_736_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_740_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_736_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_736_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_736_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_740_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_736_inst_ack_1, ack => convolution3D_CP_1120_elements(66)); -- 
    rr_1754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(66), ack => type_cast_740_inst_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_740_Sample/ra
      -- CP-element group 67: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_740_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_740_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_740_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_740_inst_ack_0, ack => convolution3D_CP_1120_elements(67)); -- 
    -- CP-element group 68:  fork  transition  place  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	64 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	201 
    -- CP-element group 68: 	202 
    -- CP-element group 68:  members (11) 
      -- CP-element group 68: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_740_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/$exit
      -- CP-element group 68: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_740_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741/type_cast_740_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_435/assign_stmt_728_to_assign_stmt_741__exit__
      -- CP-element group 68: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi
      -- CP-element group 68: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_744/$entry
      -- CP-element group 68: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_751/$entry
      -- CP-element group 68: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_740_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_740_inst_ack_1, ack => convolution3D_CP_1120_elements(68)); -- 
    -- CP-element group 69:  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	207 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/RPIPE_maxpool_input_pipe_760_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/RPIPE_maxpool_input_pipe_760_update_start_
      -- CP-element group 69: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/RPIPE_maxpool_input_pipe_760_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/RPIPE_maxpool_input_pipe_760_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/RPIPE_maxpool_input_pipe_760_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/RPIPE_maxpool_input_pipe_760_Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_760_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_760_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_1772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_760_inst_ack_0, ack => convolution3D_CP_1120_elements(69)); -- 
    cr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(69), ack => RPIPE_maxpool_input_pipe_760_inst_req_1); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/RPIPE_maxpool_input_pipe_760_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/type_cast_764_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/RPIPE_maxpool_input_pipe_760_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/RPIPE_maxpool_input_pipe_760_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/type_cast_764_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/type_cast_764_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(70) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_760_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_764_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_760_inst_ack_1, ack => convolution3D_CP_1120_elements(70)); -- 
    rr_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(70), ack => type_cast_764_inst_req_0); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/type_cast_764_Sample/ra
      -- CP-element group 71: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/type_cast_764_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/type_cast_764_Sample/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(71) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_764_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_764_inst_ack_0, ack => convolution3D_CP_1120_elements(71)); -- 
    -- CP-element group 72:  branch  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	207 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (13) 
      -- CP-element group 72: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/$exit
      -- CP-element group 72: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/type_cast_764_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/type_cast_764_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/type_cast_764_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_435/if_stmt_788_dead_link/$entry
      -- CP-element group 72: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787__exit__
      -- CP-element group 72: 	 branch_block_stmt_435/if_stmt_788__entry__
      -- CP-element group 72: 	 branch_block_stmt_435/if_stmt_788_eval_test/$entry
      -- CP-element group 72: 	 branch_block_stmt_435/if_stmt_788_eval_test/$exit
      -- CP-element group 72: 	 branch_block_stmt_435/if_stmt_788_eval_test/branch_req
      -- CP-element group 72: 	 branch_block_stmt_435/R_exitcond2_789_place
      -- CP-element group 72: 	 branch_block_stmt_435/if_stmt_788_if_link/$entry
      -- CP-element group 72: 	 branch_block_stmt_435/if_stmt_788_else_link/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(72) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_764_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_788_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_764_inst_ack_1, ack => convolution3D_CP_1120_elements(72)); -- 
    branch_req_1799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(72), ack => if_stmt_788_branch_req_0); -- 
    -- CP-element group 73:  fork  transition  place  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	208 
    -- CP-element group 73: 	209 
    -- CP-element group 73:  members (12) 
      -- CP-element group 73: 	 branch_block_stmt_435/if_stmt_788_if_link/$exit
      -- CP-element group 73: 	 branch_block_stmt_435/if_stmt_788_if_link/if_choice_transition
      -- CP-element group 73: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 73: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 73: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/$entry
      -- CP-element group 73: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/$entry
      -- CP-element group 73: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/type_cast_798/$entry
      -- CP-element group 73: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/type_cast_798/SplitProtocol/$entry
      -- CP-element group 73: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/type_cast_798/SplitProtocol/Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/type_cast_798/SplitProtocol/Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/type_cast_798/SplitProtocol/Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/type_cast_798/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_788_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_798_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_798_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_1804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_788_branch_ack_1, ack => convolution3D_CP_1120_elements(73)); -- 
    rr_2942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(73), ack => type_cast_798_inst_req_0); -- 
    cr_2947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(73), ack => type_cast_798_inst_req_1); -- 
    -- CP-element group 74:  fork  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	194 
    -- CP-element group 74: 	195 
    -- CP-element group 74: 	197 
    -- CP-element group 74: 	198 
    -- CP-element group 74:  members (20) 
      -- CP-element group 74: 	 branch_block_stmt_435/if_stmt_788_else_link/$exit
      -- CP-element group 74: 	 branch_block_stmt_435/if_stmt_788_else_link/else_choice_transition
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/$entry
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/$entry
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_747/$entry
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_747/SplitProtocol/$entry
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_747/SplitProtocol/Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_747/SplitProtocol/Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_747/SplitProtocol/Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_747/SplitProtocol/Update/cr
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/$entry
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/$entry
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/$entry
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/$entry
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_788_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_747_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_747_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_754_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_754_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_1808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_788_branch_ack_0, ack => convolution3D_CP_1120_elements(74)); -- 
    rr_2864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(74), ack => type_cast_747_inst_req_0); -- 
    cr_2869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(74), ack => type_cast_747_inst_req_1); -- 
    rr_2887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(74), ack => type_cast_754_inst_req_0); -- 
    cr_2892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(74), ack => type_cast_754_inst_req_1); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	211 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	81 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_final_index_sum_regn_sample_complete
      -- CP-element group 75: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_final_index_sum_regn_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_827_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_827_index_offset_ack_0, ack => convolution3D_CP_1120_elements(75)); -- 
    -- CP-element group 76:  transition  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	211 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (11) 
      -- CP-element group 76: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/addr_of_828_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_root_address_calculated
      -- CP-element group 76: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_offset_calculated
      -- CP-element group 76: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_final_index_sum_regn_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_final_index_sum_regn_Update/ack
      -- CP-element group 76: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_base_plus_offset/$entry
      -- CP-element group 76: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_base_plus_offset/$exit
      -- CP-element group 76: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_base_plus_offset/sum_rename_req
      -- CP-element group 76: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_base_plus_offset/sum_rename_ack
      -- CP-element group 76: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/addr_of_828_request/$entry
      -- CP-element group 76: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/addr_of_828_request/req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_827_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_828_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_827_index_offset_ack_1, ack => convolution3D_CP_1120_elements(76)); -- 
    req_1853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(76), ack => addr_of_828_final_reg_req_0); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/addr_of_828_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/addr_of_828_request/$exit
      -- CP-element group 77: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/addr_of_828_request/ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_828_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_828_final_reg_ack_0, ack => convolution3D_CP_1120_elements(77)); -- 
    -- CP-element group 78:  join  fork  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	211 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (28) 
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/addr_of_828_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/addr_of_828_complete/$exit
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/addr_of_828_complete/ack
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_base_address_calculated
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_word_address_calculated
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_root_address_calculated
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_base_address_resized
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_base_addr_resize/$entry
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_base_addr_resize/$exit
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_base_addr_resize/base_resize_req
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_base_addr_resize/base_resize_ack
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_base_plus_offset/$entry
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_base_plus_offset/$exit
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_base_plus_offset/sum_rename_req
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_base_plus_offset/sum_rename_ack
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_word_addrgen/$entry
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_word_addrgen/$exit
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_word_addrgen/root_register_req
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_word_addrgen/root_register_ack
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Sample/ptr_deref_831_Split/$entry
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Sample/ptr_deref_831_Split/$exit
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Sample/ptr_deref_831_Split/split_req
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Sample/ptr_deref_831_Split/split_ack
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Sample/word_access_start/$entry
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Sample/word_access_start/word_0/$entry
      -- CP-element group 78: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(78) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_828_final_reg_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_831_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_828_final_reg_ack_1, ack => convolution3D_CP_1120_elements(78)); -- 
    rr_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(78), ack => ptr_deref_831_store_0_req_0); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Sample/word_access_start/$exit
      -- CP-element group 79: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Sample/word_access_start/word_0/$exit
      -- CP-element group 79: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_831_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_831_store_0_ack_0, ack => convolution3D_CP_1120_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	211 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Update/word_access_complete/$exit
      -- CP-element group 80: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Update/word_access_complete/word_0/$exit
      -- CP-element group 80: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_831_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_831_store_0_ack_1, ack => convolution3D_CP_1120_elements(80)); -- 
    -- CP-element group 81:  join  transition  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	212 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833__exit__
      -- CP-element group 81: 	 branch_block_stmt_435/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 81: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/$exit
      -- CP-element group 81: 	 branch_block_stmt_435/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- CP-element group 81: 	 branch_block_stmt_435/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(81) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(75) & convolution3D_CP_1120_elements(80);
      gj_convolution3D_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	212 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_838_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_838_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_838_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_838_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_838_inst_ack_0, ack => convolution3D_CP_1120_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	212 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	88 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_838_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_838_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_838_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(83) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_838_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_838_inst_ack_1, ack => convolution3D_CP_1120_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	212 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_842_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_842_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_842_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(84) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_842_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_0, ack => convolution3D_CP_1120_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	212 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	88 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_842_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_842_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_842_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(85) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_842_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_1, ack => convolution3D_CP_1120_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	212 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_846_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_846_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_846_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(86) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_846_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_846_inst_ack_0, ack => convolution3D_CP_1120_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	212 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_846_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_846_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_846_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(87) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_846_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_846_inst_ack_1, ack => convolution3D_CP_1120_elements(87)); -- 
    -- CP-element group 88:  branch  join  transition  place  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	83 
    -- CP-element group 88: 	85 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (10) 
      -- CP-element group 88: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883__exit__
      -- CP-element group 88: 	 branch_block_stmt_435/if_stmt_884__entry__
      -- CP-element group 88: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/$exit
      -- CP-element group 88: 	 branch_block_stmt_435/if_stmt_884_dead_link/$entry
      -- CP-element group 88: 	 branch_block_stmt_435/if_stmt_884_eval_test/$entry
      -- CP-element group 88: 	 branch_block_stmt_435/if_stmt_884_eval_test/$exit
      -- CP-element group 88: 	 branch_block_stmt_435/if_stmt_884_eval_test/branch_req
      -- CP-element group 88: 	 branch_block_stmt_435/R_cmp65191_885_place
      -- CP-element group 88: 	 branch_block_stmt_435/if_stmt_884_if_link/$entry
      -- CP-element group 88: 	 branch_block_stmt_435/if_stmt_884_else_link/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_884_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(88), ack => if_stmt_884_branch_req_0); -- 
    convolution3D_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(83) & convolution3D_CP_1120_elements(85) & convolution3D_CP_1120_elements(87);
      gj_convolution3D_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: 	92 
    -- CP-element group 89: 	93 
    -- CP-element group 89: 	94 
    -- CP-element group 89: 	95 
    -- CP-element group 89: 	96 
    -- CP-element group 89: 	97 
    -- CP-element group 89: 	98 
    -- CP-element group 89: 	101 
    -- CP-element group 89: 	103 
    -- CP-element group 89:  members (42) 
      -- CP-element group 89: 	 branch_block_stmt_435/merge_stmt_890__exit__
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961__entry__
      -- CP-element group 89: 	 branch_block_stmt_435/if_stmt_884_if_link/$exit
      -- CP-element group 89: 	 branch_block_stmt_435/if_stmt_884_if_link/if_choice_transition
      -- CP-element group 89: 	 branch_block_stmt_435/ifx_xend_bbx_xnph
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/$entry
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_905_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_905_update_start_
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_905_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_905_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_905_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_905_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_909_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_909_update_start_
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_909_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_909_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_909_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_909_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_918_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_918_update_start_
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_918_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_918_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_918_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_918_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_927_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_927_update_start_
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_927_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_927_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_927_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_927_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_936_update_start_
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_936_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_936_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_941_update_start_
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_941_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_941_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_435/ifx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 89: 	 branch_block_stmt_435/ifx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 89: 	 branch_block_stmt_435/merge_stmt_890_PhiReqMerge
      -- CP-element group 89: 	 branch_block_stmt_435/merge_stmt_890_PhiAck/$entry
      -- CP-element group 89: 	 branch_block_stmt_435/merge_stmt_890_PhiAck/$exit
      -- CP-element group 89: 	 branch_block_stmt_435/merge_stmt_890_PhiAck/dummy
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_884_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_905_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_905_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_909_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_909_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_918_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_918_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_927_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_927_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_936_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_941_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_1967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_884_branch_ack_1, ack => convolution3D_CP_1120_elements(89)); -- 
    rr_1984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(89), ack => type_cast_905_inst_req_0); -- 
    cr_1989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(89), ack => type_cast_905_inst_req_1); -- 
    rr_1998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(89), ack => type_cast_909_inst_req_0); -- 
    cr_2003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(89), ack => type_cast_909_inst_req_1); -- 
    rr_2012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(89), ack => type_cast_918_inst_req_0); -- 
    cr_2017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(89), ack => type_cast_918_inst_req_1); -- 
    rr_2026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(89), ack => type_cast_927_inst_req_0); -- 
    cr_2031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(89), ack => type_cast_927_inst_req_1); -- 
    cr_2045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(89), ack => type_cast_936_inst_req_1); -- 
    cr_2059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(89), ack => type_cast_941_inst_req_1); -- 
    -- CP-element group 90:  transition  place  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	222 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_435/if_stmt_884_else_link/$exit
      -- CP-element group 90: 	 branch_block_stmt_435/if_stmt_884_else_link/else_choice_transition
      -- CP-element group 90: 	 branch_block_stmt_435/ifx_xend_forx_xend95
      -- CP-element group 90: 	 branch_block_stmt_435/ifx_xend_forx_xend95_PhiReq/$entry
      -- CP-element group 90: 	 branch_block_stmt_435/ifx_xend_forx_xend95_PhiReq/phi_stmt_1086/$entry
      -- CP-element group 90: 	 branch_block_stmt_435/ifx_xend_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(90) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_884_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_1971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_884_branch_ack_0, ack => convolution3D_CP_1120_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_905_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_905_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_905_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(91) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_905_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_0, ack => convolution3D_CP_1120_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	89 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	99 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_905_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_905_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_905_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(92) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_905_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_1, ack => convolution3D_CP_1120_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	89 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_909_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_909_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_909_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_909_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_909_inst_ack_0, ack => convolution3D_CP_1120_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	89 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	99 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_909_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_909_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_909_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_909_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_909_inst_ack_1, ack => convolution3D_CP_1120_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	89 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_918_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_918_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_918_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(95) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_918_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_918_inst_ack_0, ack => convolution3D_CP_1120_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	89 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	99 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_918_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_918_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_918_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(96) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_918_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_918_inst_ack_1, ack => convolution3D_CP_1120_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	89 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_927_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_927_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_927_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(97) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_927_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_0, ack => convolution3D_CP_1120_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	89 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_927_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_927_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_927_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_927_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_1, ack => convolution3D_CP_1120_elements(98)); -- 
    -- CP-element group 99:  join  transition  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	92 
    -- CP-element group 99: 	94 
    -- CP-element group 99: 	96 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_936_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_936_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_936_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(99) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_936_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(99), ack => type_cast_936_inst_req_0); -- 
    convolution3D_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(92) & convolution3D_CP_1120_elements(94) & convolution3D_CP_1120_elements(96) & convolution3D_CP_1120_elements(98);
      gj_convolution3D_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_936_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_936_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_936_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(100) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_936_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_936_inst_ack_0, ack => convolution3D_CP_1120_elements(100)); -- 
    -- CP-element group 101:  transition  input  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	89 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (6) 
      -- CP-element group 101: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_936_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_936_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_936_Update/ca
      -- CP-element group 101: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_941_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_941_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_941_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(101) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_936_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_941_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_2046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_936_inst_ack_1, ack => convolution3D_CP_1120_elements(101)); -- 
    rr_2054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(101), ack => type_cast_941_inst_req_0); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_941_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_941_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_941_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(102) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_941_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_941_inst_ack_0, ack => convolution3D_CP_1120_elements(102)); -- 
    -- CP-element group 103:  transition  place  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	89 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	213 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961__exit__
      -- CP-element group 103: 	 branch_block_stmt_435/bbx_xnph_forx_xbody67
      -- CP-element group 103: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/$exit
      -- CP-element group 103: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_941_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_941_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_435/assign_stmt_896_to_assign_stmt_961/type_cast_941_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_435/bbx_xnph_forx_xbody67_PhiReq/$entry
      -- CP-element group 103: 	 branch_block_stmt_435/bbx_xnph_forx_xbody67_PhiReq/phi_stmt_964/$entry
      -- CP-element group 103: 	 branch_block_stmt_435/bbx_xnph_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(103) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_941_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_941_inst_ack_1, ack => convolution3D_CP_1120_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	218 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	127 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_final_index_sum_regn_sample_complete
      -- CP-element group 104: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_final_index_sum_regn_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(104) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_976_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_976_index_offset_ack_0, ack => convolution3D_CP_1120_elements(104)); -- 
    -- CP-element group 105:  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	218 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (11) 
      -- CP-element group 105: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/addr_of_977_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_root_address_calculated
      -- CP-element group 105: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_offset_calculated
      -- CP-element group 105: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_final_index_sum_regn_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_final_index_sum_regn_Update/ack
      -- CP-element group 105: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_base_plus_offset/$entry
      -- CP-element group 105: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_base_plus_offset/$exit
      -- CP-element group 105: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_base_plus_offset/sum_rename_req
      -- CP-element group 105: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_base_plus_offset/sum_rename_ack
      -- CP-element group 105: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/addr_of_977_request/$entry
      -- CP-element group 105: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/addr_of_977_request/req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(105) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_976_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_977_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_976_index_offset_ack_1, ack => convolution3D_CP_1120_elements(105)); -- 
    req_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(105), ack => addr_of_977_final_reg_req_0); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/addr_of_977_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/addr_of_977_request/$exit
      -- CP-element group 106: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/addr_of_977_request/ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(106) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_977_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_977_final_reg_ack_0, ack => convolution3D_CP_1120_elements(106)); -- 
    -- CP-element group 107:  fork  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	218 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	124 
    -- CP-element group 107:  members (19) 
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/addr_of_977_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/addr_of_977_complete/$exit
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/addr_of_977_complete/ack
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_base_address_calculated
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_word_address_calculated
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_root_address_calculated
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_base_address_resized
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_base_addr_resize/$entry
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_base_addr_resize/$exit
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_base_addr_resize/base_resize_req
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_base_addr_resize/base_resize_ack
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_base_plus_offset/$entry
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_base_plus_offset/$exit
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_base_plus_offset/sum_rename_req
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_base_plus_offset/sum_rename_ack
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_word_addrgen/$entry
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_word_addrgen/$exit
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_word_addrgen/root_register_req
      -- CP-element group 107: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(107)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(107)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(107) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_977_final_reg_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_977_final_reg_ack_1, ack => convolution3D_CP_1120_elements(107)); -- 
    -- CP-element group 108:  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	218 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (6) 
      -- CP-element group 108: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_980_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_980_update_start_
      -- CP-element group 108: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_980_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_980_Sample/ra
      -- CP-element group 108: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_980_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_980_Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(108)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(108)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(108) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_980_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_980_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_2118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_980_inst_ack_0, ack => convolution3D_CP_1120_elements(108)); -- 
    cr_2122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(108), ack => RPIPE_maxpool_input_pipe_980_inst_req_1); -- 
    -- CP-element group 109:  fork  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: 	112 
    -- CP-element group 109:  members (9) 
      -- CP-element group 109: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_980_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_980_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_980_Update/ca
      -- CP-element group 109: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_984_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_984_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_984_Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_993_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_993_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_993_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(109)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(109)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(109) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_980_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_984_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_993_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_2123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_980_inst_ack_1, ack => convolution3D_CP_1120_elements(109)); -- 
    rr_2131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(109), ack => type_cast_984_inst_req_0); -- 
    rr_2145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(109), ack => RPIPE_maxpool_input_pipe_993_inst_req_0); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_984_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_984_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_984_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(110)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(110)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(110) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_984_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_984_inst_ack_0, ack => convolution3D_CP_1120_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	218 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	124 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_984_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_984_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_984_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(111)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(111)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(111) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_984_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_984_inst_ack_1, ack => convolution3D_CP_1120_elements(111)); -- 
    -- CP-element group 112:  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	109 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (6) 
      -- CP-element group 112: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_993_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_993_update_start_
      -- CP-element group 112: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_993_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_993_Sample/ra
      -- CP-element group 112: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_993_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_993_Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(112)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(112)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(112) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_993_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_993_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_2146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_993_inst_ack_0, ack => convolution3D_CP_1120_elements(112)); -- 
    cr_2150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(112), ack => RPIPE_maxpool_input_pipe_993_inst_req_1); -- 
    -- CP-element group 113:  fork  transition  input  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113: 	116 
    -- CP-element group 113:  members (9) 
      -- CP-element group 113: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_993_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_993_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_993_Update/ca
      -- CP-element group 113: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_997_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_997_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_997_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1011_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1011_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1011_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(113)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(113)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(113) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_993_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_997_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_1011_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_2151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_993_inst_ack_1, ack => convolution3D_CP_1120_elements(113)); -- 
    rr_2159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(113), ack => type_cast_997_inst_req_0); -- 
    rr_2173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(113), ack => RPIPE_maxpool_input_pipe_1011_inst_req_0); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_997_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_997_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_997_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(114)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(114)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(114) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_997_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_997_inst_ack_0, ack => convolution3D_CP_1120_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	218 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	124 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_997_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_997_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_997_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(115)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(115)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(115) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_997_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_997_inst_ack_1, ack => convolution3D_CP_1120_elements(115)); -- 
    -- CP-element group 116:  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	113 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (6) 
      -- CP-element group 116: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1011_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1011_update_start_
      -- CP-element group 116: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1011_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1011_Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1011_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1011_Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(116)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(116)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(116) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_1011_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_1011_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_2174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1011_inst_ack_0, ack => convolution3D_CP_1120_elements(116)); -- 
    cr_2178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(116), ack => RPIPE_maxpool_input_pipe_1011_inst_req_1); -- 
    -- CP-element group 117:  fork  transition  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117: 	120 
    -- CP-element group 117:  members (9) 
      -- CP-element group 117: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1011_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1011_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1011_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1015_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1015_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1015_Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1029_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1029_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1029_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(117)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(117)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(117) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_1011_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1015_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_1029_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_2179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1011_inst_ack_1, ack => convolution3D_CP_1120_elements(117)); -- 
    rr_2187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(117), ack => type_cast_1015_inst_req_0); -- 
    rr_2201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(117), ack => RPIPE_maxpool_input_pipe_1029_inst_req_0); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1015_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1015_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1015_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(118)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(118)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(118) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1015_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1015_inst_ack_0, ack => convolution3D_CP_1120_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	218 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1015_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1015_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1015_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(119)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(119)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(119) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1015_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1015_inst_ack_1, ack => convolution3D_CP_1120_elements(119)); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	117 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1029_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1029_update_start_
      -- CP-element group 120: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1029_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1029_Sample/ra
      -- CP-element group 120: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1029_Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1029_Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(120)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(120)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(120) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_1029_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_1029_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_2202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1029_inst_ack_0, ack => convolution3D_CP_1120_elements(120)); -- 
    cr_2206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(120), ack => RPIPE_maxpool_input_pipe_1029_inst_req_1); -- 
    -- CP-element group 121:  transition  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (6) 
      -- CP-element group 121: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1029_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1029_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_1029_Update/ca
      -- CP-element group 121: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1033_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1033_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1033_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(121)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(121)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(121) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_1029_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1033_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_2207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1029_inst_ack_1, ack => convolution3D_CP_1120_elements(121)); -- 
    rr_2215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(121), ack => type_cast_1033_inst_req_0); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1033_sample_completed_
      -- CP-element group 122: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1033_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1033_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(122)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(122)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(122) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1033_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1033_inst_ack_0, ack => convolution3D_CP_1120_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	218 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1033_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1033_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1033_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(123)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(123)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(123) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1033_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1033_inst_ack_1, ack => convolution3D_CP_1120_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	107 
    -- CP-element group 124: 	111 
    -- CP-element group 124: 	115 
    -- CP-element group 124: 	119 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Sample/ptr_deref_1041_Split/$entry
      -- CP-element group 124: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Sample/ptr_deref_1041_Split/$exit
      -- CP-element group 124: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Sample/ptr_deref_1041_Split/split_req
      -- CP-element group 124: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Sample/ptr_deref_1041_Split/split_ack
      -- CP-element group 124: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Sample/word_access_start/$entry
      -- CP-element group 124: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Sample/word_access_start/word_0/$entry
      -- CP-element group 124: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(124)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(124)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(124) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_1041_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(124), ack => ptr_deref_1041_store_0_req_0); -- 
    convolution3D_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(107) & convolution3D_CP_1120_elements(111) & convolution3D_CP_1120_elements(115) & convolution3D_CP_1120_elements(119) & convolution3D_CP_1120_elements(123);
      gj_convolution3D_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Sample/word_access_start/$exit
      -- CP-element group 125: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Sample/word_access_start/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(125)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(125)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(125) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_1041_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_store_0_ack_0, ack => convolution3D_CP_1120_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	218 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Update/word_access_complete/$exit
      -- CP-element group 126: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Update/word_access_complete/word_0/$exit
      -- CP-element group 126: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(126)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(126)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(126) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_1041_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_store_0_ack_1, ack => convolution3D_CP_1120_elements(126)); -- 
    -- CP-element group 127:  branch  join  transition  place  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	104 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (10) 
      -- CP-element group 127: 	 branch_block_stmt_435/if_stmt_1055_eval_test/branch_req
      -- CP-element group 127: 	 branch_block_stmt_435/if_stmt_1055_eval_test/$exit
      -- CP-element group 127: 	 branch_block_stmt_435/if_stmt_1055_if_link/$entry
      -- CP-element group 127: 	 branch_block_stmt_435/if_stmt_1055_eval_test/$entry
      -- CP-element group 127: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054__exit__
      -- CP-element group 127: 	 branch_block_stmt_435/if_stmt_1055__entry__
      -- CP-element group 127: 	 branch_block_stmt_435/R_exitcond26_1056_place
      -- CP-element group 127: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/$exit
      -- CP-element group 127: 	 branch_block_stmt_435/if_stmt_1055_else_link/$entry
      -- CP-element group 127: 	 branch_block_stmt_435/if_stmt_1055_dead_link/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(127)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(127)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(127) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_1055_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_2279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(127), ack => if_stmt_1055_branch_req_0); -- 
    convolution3D_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(104) & convolution3D_CP_1120_elements(126);
      gj_convolution3D_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	219 
    -- CP-element group 128: 	220 
    -- CP-element group 128:  members (24) 
      -- CP-element group 128: 	 branch_block_stmt_435/if_stmt_1055_if_link/$exit
      -- CP-element group 128: 	 branch_block_stmt_435/merge_stmt_1061__exit__
      -- CP-element group 128: 	 branch_block_stmt_435/assign_stmt_1068_to_assign_stmt_1083__entry__
      -- CP-element group 128: 	 branch_block_stmt_435/assign_stmt_1068_to_assign_stmt_1083__exit__
      -- CP-element group 128: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95
      -- CP-element group 128: 	 branch_block_stmt_435/if_stmt_1055_if_link/if_choice_transition
      -- CP-element group 128: 	 branch_block_stmt_435/assign_stmt_1068_to_assign_stmt_1083/$exit
      -- CP-element group 128: 	 branch_block_stmt_435/forx_xbody67_forx_xcond60x_xforx_xend95_crit_edge
      -- CP-element group 128: 	 branch_block_stmt_435/assign_stmt_1068_to_assign_stmt_1083/$entry
      -- CP-element group 128: 	 branch_block_stmt_435/forx_xbody67_forx_xcond60x_xforx_xend95_crit_edge_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_435/forx_xbody67_forx_xcond60x_xforx_xend95_crit_edge_PhiReq/$exit
      -- CP-element group 128: 	 branch_block_stmt_435/merge_stmt_1061_PhiReqMerge
      -- CP-element group 128: 	 branch_block_stmt_435/merge_stmt_1061_PhiAck/$entry
      -- CP-element group 128: 	 branch_block_stmt_435/merge_stmt_1061_PhiAck/$exit
      -- CP-element group 128: 	 branch_block_stmt_435/merge_stmt_1061_PhiAck/dummy
      -- CP-element group 128: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/$entry
      -- CP-element group 128: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/type_cast_1089/$entry
      -- CP-element group 128: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/type_cast_1089/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/type_cast_1089/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/type_cast_1089/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/type_cast_1089/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/type_cast_1089/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(128)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(128)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(128) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_1055_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1089_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1089_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_2284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1055_branch_ack_1, ack => convolution3D_CP_1120_elements(128)); -- 
    rr_3050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(128), ack => type_cast_1089_inst_req_0); -- 
    cr_3055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(128), ack => type_cast_1089_inst_req_1); -- 
    -- CP-element group 129:  fork  transition  place  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	214 
    -- CP-element group 129: 	215 
    -- CP-element group 129:  members (12) 
      -- CP-element group 129: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67
      -- CP-element group 129: 	 branch_block_stmt_435/if_stmt_1055_else_link/else_choice_transition
      -- CP-element group 129: 	 branch_block_stmt_435/if_stmt_1055_else_link/$exit
      -- CP-element group 129: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/$entry
      -- CP-element group 129: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/$entry
      -- CP-element group 129: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/$entry
      -- CP-element group 129: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/type_cast_970/$entry
      -- CP-element group 129: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/type_cast_970/SplitProtocol/$entry
      -- CP-element group 129: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/type_cast_970/SplitProtocol/Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/type_cast_970/SplitProtocol/Sample/rr
      -- CP-element group 129: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/type_cast_970/SplitProtocol/Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/type_cast_970/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(129)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(129)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(129) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_1055_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_970_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_970_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_2288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1055_branch_ack_0, ack => convolution3D_CP_1120_elements(129)); -- 
    rr_3007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(129), ack => type_cast_970_inst_req_0); -- 
    cr_3012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(129), ack => type_cast_970_inst_req_1); -- 
    -- CP-element group 130:  transition  place  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	224 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	243 
    -- CP-element group 130:  members (5) 
      -- CP-element group 130: 	 branch_block_stmt_435/if_stmt_1106_if_link/if_choice_transition
      -- CP-element group 130: 	 branch_block_stmt_435/if_stmt_1106_if_link/$exit
      -- CP-element group 130: 	 branch_block_stmt_435/forx_xend95_ifx_xend107
      -- CP-element group 130: 	 branch_block_stmt_435/forx_xend95_ifx_xend107_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_435/forx_xend95_ifx_xend107_PhiReq/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(130)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(130)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(130) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_1106_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_2309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1106_branch_ack_1, ack => convolution3D_CP_1120_elements(130)); -- 
    -- CP-element group 131:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	224 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131: 	133 
    -- CP-element group 131: 	135 
    -- CP-element group 131:  members (21) 
      -- CP-element group 131: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1130_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1134_update_start_
      -- CP-element group 131: 	 branch_block_stmt_435/if_stmt_1106_else_link/$exit
      -- CP-element group 131: 	 branch_block_stmt_435/if_stmt_1106_else_link/else_choice_transition
      -- CP-element group 131: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/$entry
      -- CP-element group 131: 	 branch_block_stmt_435/merge_stmt_1112__exit__
      -- CP-element group 131: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1130_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135__entry__
      -- CP-element group 131: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1130_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_435/forx_xend95_forx_xbodyx_xi181x_xpreheader
      -- CP-element group 131: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1134_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1130_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1130_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1130_update_start_
      -- CP-element group 131: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1134_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_435/forx_xend95_forx_xbodyx_xi181x_xpreheader_PhiReq/$entry
      -- CP-element group 131: 	 branch_block_stmt_435/forx_xend95_forx_xbodyx_xi181x_xpreheader_PhiReq/$exit
      -- CP-element group 131: 	 branch_block_stmt_435/merge_stmt_1112_PhiReqMerge
      -- CP-element group 131: 	 branch_block_stmt_435/merge_stmt_1112_PhiAck/$entry
      -- CP-element group 131: 	 branch_block_stmt_435/merge_stmt_1112_PhiAck/$exit
      -- CP-element group 131: 	 branch_block_stmt_435/merge_stmt_1112_PhiAck/dummy
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(131)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(131)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(131) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_1106_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1130_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1134_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1130_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_2313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1106_branch_ack_0, ack => convolution3D_CP_1120_elements(131)); -- 
    cr_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(131), ack => type_cast_1130_inst_req_1); -- 
    cr_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(131), ack => type_cast_1134_inst_req_1); -- 
    rr_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(131), ack => type_cast_1130_inst_req_0); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1130_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1130_Sample/ra
      -- CP-element group 132: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1130_Sample/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(132)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(132)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(132) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1130_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1130_inst_ack_0, ack => convolution3D_CP_1120_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1134_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1130_Update/ca
      -- CP-element group 133: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1134_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1130_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1130_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1134_Sample/rr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(133)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(133)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(133) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1130_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1134_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1130_inst_ack_1, ack => convolution3D_CP_1120_elements(133)); -- 
    rr_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(133), ack => type_cast_1134_inst_req_0); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1134_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1134_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1134_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(134)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(134)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(134) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1134_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1134_inst_ack_0, ack => convolution3D_CP_1120_elements(134)); -- 
    -- CP-element group 135:  fork  transition  place  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	131 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	232 
    -- CP-element group 135: 	233 
    -- CP-element group 135:  members (11) 
      -- CP-element group 135: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/$exit
      -- CP-element group 135: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135__exit__
      -- CP-element group 135: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181
      -- CP-element group 135: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1134_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1134_Update/ca
      -- CP-element group 135: 	 branch_block_stmt_435/assign_stmt_1117_to_assign_stmt_1135/type_cast_1134_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/$entry
      -- CP-element group 135: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/$entry
      -- CP-element group 135: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/$entry
      -- CP-element group 135: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/$entry
      -- CP-element group 135: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(135)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(135)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(135) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1134_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1134_inst_ack_1, ack => convolution3D_CP_1120_elements(135)); -- 
    -- CP-element group 136:  transition  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	238 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (6) 
      -- CP-element group 136: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/RPIPE_maxpool_input_pipe_1154_update_start_
      -- CP-element group 136: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/RPIPE_maxpool_input_pipe_1154_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/RPIPE_maxpool_input_pipe_1154_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/RPIPE_maxpool_input_pipe_1154_Update/cr
      -- CP-element group 136: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/RPIPE_maxpool_input_pipe_1154_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/RPIPE_maxpool_input_pipe_1154_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(136)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(136)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(136) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_1154_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_1154_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_2358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1154_inst_ack_0, ack => convolution3D_CP_1120_elements(136)); -- 
    cr_2362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(136), ack => RPIPE_maxpool_input_pipe_1154_inst_req_1); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/RPIPE_maxpool_input_pipe_1154_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/type_cast_1158_Sample/rr
      -- CP-element group 137: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/type_cast_1158_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/type_cast_1158_sample_start_
      -- CP-element group 137: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/RPIPE_maxpool_input_pipe_1154_Update/ca
      -- CP-element group 137: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/RPIPE_maxpool_input_pipe_1154_Update/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(137)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(137)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(137) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_1154_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1158_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_2363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1154_inst_ack_1, ack => convolution3D_CP_1120_elements(137)); -- 
    rr_2371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(137), ack => type_cast_1158_inst_req_0); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/type_cast_1158_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/type_cast_1158_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/type_cast_1158_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(138)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(138)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(138) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1158_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1158_inst_ack_0, ack => convolution3D_CP_1120_elements(138)); -- 
    -- CP-element group 139:  branch  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	238 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (13) 
      -- CP-element group 139: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181__exit__
      -- CP-element group 139: 	 branch_block_stmt_435/if_stmt_1182__entry__
      -- CP-element group 139: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/$exit
      -- CP-element group 139: 	 branch_block_stmt_435/if_stmt_1182_else_link/$entry
      -- CP-element group 139: 	 branch_block_stmt_435/R_exitcond_1183_place
      -- CP-element group 139: 	 branch_block_stmt_435/if_stmt_1182_if_link/$entry
      -- CP-element group 139: 	 branch_block_stmt_435/if_stmt_1182_eval_test/branch_req
      -- CP-element group 139: 	 branch_block_stmt_435/if_stmt_1182_eval_test/$exit
      -- CP-element group 139: 	 branch_block_stmt_435/if_stmt_1182_eval_test/$entry
      -- CP-element group 139: 	 branch_block_stmt_435/if_stmt_1182_dead_link/$entry
      -- CP-element group 139: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/type_cast_1158_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/type_cast_1158_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/type_cast_1158_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(139)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(139)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(139) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1158_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_1182_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_2377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1158_inst_ack_1, ack => convolution3D_CP_1120_elements(139)); -- 
    branch_req_2385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(139), ack => if_stmt_1182_branch_req_0); -- 
    -- CP-element group 140:  fork  transition  place  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	239 
    -- CP-element group 140: 	240 
    -- CP-element group 140:  members (12) 
      -- CP-element group 140: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188
      -- CP-element group 140: 	 branch_block_stmt_435/if_stmt_1182_if_link/if_choice_transition
      -- CP-element group 140: 	 branch_block_stmt_435/if_stmt_1182_if_link/$exit
      -- CP-element group 140: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/$entry
      -- CP-element group 140: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/$entry
      -- CP-element group 140: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/$entry
      -- CP-element group 140: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/type_cast_1192/$entry
      -- CP-element group 140: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/type_cast_1192/SplitProtocol/$entry
      -- CP-element group 140: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/type_cast_1192/SplitProtocol/Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/type_cast_1192/SplitProtocol/Sample/rr
      -- CP-element group 140: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/type_cast_1192/SplitProtocol/Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/type_cast_1192/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(140)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(140)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(140) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_1182_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1192_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1192_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_2390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1182_branch_ack_1, ack => convolution3D_CP_1120_elements(140)); -- 
    rr_3182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(140), ack => type_cast_1192_inst_req_0); -- 
    cr_3187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(140), ack => type_cast_1192_inst_req_1); -- 
    -- CP-element group 141:  fork  transition  place  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	225 
    -- CP-element group 141: 	226 
    -- CP-element group 141: 	228 
    -- CP-element group 141: 	229 
    -- CP-element group 141:  members (20) 
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181
      -- CP-element group 141: 	 branch_block_stmt_435/if_stmt_1182_else_link/else_choice_transition
      -- CP-element group 141: 	 branch_block_stmt_435/if_stmt_1182_else_link/$exit
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/$entry
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/$entry
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/$entry
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/type_cast_1141/$entry
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/type_cast_1141/SplitProtocol/$entry
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/type_cast_1141/SplitProtocol/Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/type_cast_1141/SplitProtocol/Sample/rr
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/type_cast_1141/SplitProtocol/Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/type_cast_1141/SplitProtocol/Update/cr
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/$entry
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/$entry
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/type_cast_1148/$entry
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/type_cast_1148/SplitProtocol/$entry
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/type_cast_1148/SplitProtocol/Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/type_cast_1148/SplitProtocol/Sample/rr
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/type_cast_1148/SplitProtocol/Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/type_cast_1148/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(141)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(141)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(141) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_1182_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1141_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1141_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1148_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1148_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_2394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1182_branch_ack_0, ack => convolution3D_CP_1120_elements(141)); -- 
    rr_3104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(141), ack => type_cast_1141_inst_req_0); -- 
    cr_3109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(141), ack => type_cast_1141_inst_req_1); -- 
    rr_3127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(141), ack => type_cast_1148_inst_req_0); -- 
    cr_3132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(141), ack => type_cast_1148_inst_req_1); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	242 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	148 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_final_index_sum_regn_Sample/ack
      -- CP-element group 142: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_final_index_sum_regn_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_final_index_sum_regn_sample_complete
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(142)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(142)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(142) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_1221_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1221_index_offset_ack_0, ack => convolution3D_CP_1120_elements(142)); -- 
    -- CP-element group 143:  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	242 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (11) 
      -- CP-element group 143: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/addr_of_1222_request/$entry
      -- CP-element group 143: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_base_plus_offset/sum_rename_ack
      -- CP-element group 143: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/addr_of_1222_request/req
      -- CP-element group 143: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_base_plus_offset/sum_rename_req
      -- CP-element group 143: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_base_plus_offset/$exit
      -- CP-element group 143: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_base_plus_offset/$entry
      -- CP-element group 143: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_offset_calculated
      -- CP-element group 143: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_final_index_sum_regn_Update/ack
      -- CP-element group 143: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_root_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/addr_of_1222_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_final_index_sum_regn_Update/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(143)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(143)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(143) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_1221_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_1222_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1221_index_offset_ack_1, ack => convolution3D_CP_1120_elements(143)); -- 
    req_2439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(143), ack => addr_of_1222_final_reg_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/addr_of_1222_request/$exit
      -- CP-element group 144: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/addr_of_1222_request/ack
      -- CP-element group 144: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/addr_of_1222_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(144)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(144)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(144) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_1222_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1222_final_reg_ack_0, ack => convolution3D_CP_1120_elements(144)); -- 
    -- CP-element group 145:  join  fork  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	242 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (28) 
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/addr_of_1222_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Sample/word_access_start/word_0/rr
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Sample/word_access_start/word_0/$entry
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Sample/word_access_start/$entry
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Sample/ptr_deref_1225_Split/split_ack
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Sample/ptr_deref_1225_Split/split_req
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Sample/ptr_deref_1225_Split/$exit
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Sample/ptr_deref_1225_Split/$entry
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_word_addrgen/root_register_ack
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_word_addrgen/root_register_req
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_word_addrgen/$exit
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_word_addrgen/$entry
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_base_plus_offset/sum_rename_ack
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_base_plus_offset/sum_rename_req
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_base_plus_offset/$exit
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_base_plus_offset/$entry
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_base_addr_resize/base_resize_ack
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_base_addr_resize/base_resize_req
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_base_addr_resize/$exit
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_base_addr_resize/$entry
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_base_address_resized
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_root_address_calculated
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_word_address_calculated
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_base_address_calculated
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/addr_of_1222_complete/ack
      -- CP-element group 145: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/addr_of_1222_complete/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(145)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(145)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(145) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_1222_final_reg_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_1225_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1222_final_reg_ack_1, ack => convolution3D_CP_1120_elements(145)); -- 
    rr_2483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(145), ack => ptr_deref_1225_store_0_req_0); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Sample/word_access_start/word_0/ra
      -- CP-element group 146: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Sample/word_access_start/word_0/$exit
      -- CP-element group 146: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Sample/word_access_start/$exit
      -- CP-element group 146: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(146)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(146)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(146) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_1225_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1225_store_0_ack_0, ack => convolution3D_CP_1120_elements(146)); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	242 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Update/word_access_complete/word_0/ca
      -- CP-element group 147: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Update/word_access_complete/word_0/$exit
      -- CP-element group 147: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Update/word_access_complete/$exit
      -- CP-element group 147: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(147)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(147)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(147) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_1225_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1225_store_0_ack_1, ack => convolution3D_CP_1120_elements(147)); -- 
    -- CP-element group 148:  join  transition  place  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	142 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	243 
    -- CP-element group 148:  members (5) 
      -- CP-element group 148: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227__exit__
      -- CP-element group 148: 	 branch_block_stmt_435/getRemainingElementsx_xexit188_ifx_xend107
      -- CP-element group 148: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/$exit
      -- CP-element group 148: 	 branch_block_stmt_435/getRemainingElementsx_xexit188_ifx_xend107_PhiReq/$entry
      -- CP-element group 148: 	 branch_block_stmt_435/getRemainingElementsx_xexit188_ifx_xend107_PhiReq/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(148)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(148)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(148) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(142) & convolution3D_CP_1120_elements(147);
      gj_convolution3D_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	243 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_435/call_stmt_1232/call_stmt_1232_Sample/cra
      -- CP-element group 149: 	 branch_block_stmt_435/call_stmt_1232/call_stmt_1232_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_435/call_stmt_1232/call_stmt_1232_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(149)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(149)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(149) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1232_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_2507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1232_call_ack_0, ack => convolution3D_CP_1120_elements(149)); -- 
    -- CP-element group 150:  fork  transition  place  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	243 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150: 	155 
    -- CP-element group 150: 	156 
    -- CP-element group 150: 	157 
    -- CP-element group 150: 	158 
    -- CP-element group 150: 	159 
    -- CP-element group 150: 	160 
    -- CP-element group 150:  members (31) 
      -- CP-element group 150: 	 branch_block_stmt_435/call_stmt_1232/call_stmt_1232_Update/cca
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/$entry
      -- CP-element group 150: 	 branch_block_stmt_435/call_stmt_1232__exit__
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296__entry__
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_num_out_pipe_1244_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_435/call_stmt_1232/call_stmt_1232_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_435/call_stmt_1232/call_stmt_1232_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1290_Update/cr
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1290_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1290_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1290_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_435/call_stmt_1232/$exit
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1290_update_start_
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1290_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1281_Update/cr
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1281_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1281_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1281_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1281_update_start_
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1281_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1271_Update/cr
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1271_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1271_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1271_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1271_update_start_
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1271_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_maxpool_output_pipe_1247_Sample/req
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_maxpool_output_pipe_1247_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_maxpool_output_pipe_1247_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_num_out_pipe_1244_Sample/req
      -- CP-element group 150: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_num_out_pipe_1244_Sample/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(150)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(150)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(150) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1232_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1290_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1290_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1281_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1281_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1271_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1271_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:WPIPE_maxpool_output_pipe_1247_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:WPIPE_num_out_pipe_1244_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_2512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1232_call_ack_1, ack => convolution3D_CP_1120_elements(150)); -- 
    cr_2584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(150), ack => type_cast_1290_inst_req_1); -- 
    rr_2579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(150), ack => type_cast_1290_inst_req_0); -- 
    cr_2570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(150), ack => type_cast_1281_inst_req_1); -- 
    rr_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(150), ack => type_cast_1281_inst_req_0); -- 
    cr_2556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(150), ack => type_cast_1271_inst_req_1); -- 
    rr_2551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(150), ack => type_cast_1271_inst_req_0); -- 
    req_2537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(150), ack => WPIPE_maxpool_output_pipe_1247_inst_req_0); -- 
    req_2523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(150), ack => WPIPE_num_out_pipe_1244_inst_req_0); -- 
    -- CP-element group 151:  transition  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151:  members (6) 
      -- CP-element group 151: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_num_out_pipe_1244_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_num_out_pipe_1244_update_start_
      -- CP-element group 151: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_num_out_pipe_1244_Update/req
      -- CP-element group 151: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_num_out_pipe_1244_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_num_out_pipe_1244_Sample/ack
      -- CP-element group 151: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_num_out_pipe_1244_Sample/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(151)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(151)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(151) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:WPIPE_num_out_pipe_1244_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:WPIPE_num_out_pipe_1244_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1244_inst_ack_0, ack => convolution3D_CP_1120_elements(151)); -- 
    req_2528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(151), ack => WPIPE_num_out_pipe_1244_inst_req_1); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_num_out_pipe_1244_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_num_out_pipe_1244_Update/ack
      -- CP-element group 152: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_num_out_pipe_1244_Update/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(152)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(152)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(152) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:WPIPE_num_out_pipe_1244_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1244_inst_ack_1, ack => convolution3D_CP_1120_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_maxpool_output_pipe_1247_Update/req
      -- CP-element group 153: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_maxpool_output_pipe_1247_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_maxpool_output_pipe_1247_Sample/ack
      -- CP-element group 153: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_maxpool_output_pipe_1247_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_maxpool_output_pipe_1247_update_start_
      -- CP-element group 153: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_maxpool_output_pipe_1247_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(153)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(153)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(153) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:WPIPE_maxpool_output_pipe_1247_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:WPIPE_maxpool_output_pipe_1247_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1247_inst_ack_0, ack => convolution3D_CP_1120_elements(153)); -- 
    req_2542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(153), ack => WPIPE_maxpool_output_pipe_1247_inst_req_1); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	161 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_maxpool_output_pipe_1247_Update/ack
      -- CP-element group 154: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_maxpool_output_pipe_1247_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/WPIPE_maxpool_output_pipe_1247_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(154)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(154)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(154) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:WPIPE_maxpool_output_pipe_1247_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1247_inst_ack_1, ack => convolution3D_CP_1120_elements(154)); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	150 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1271_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1271_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1271_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(155)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(155)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(155) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1271_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1271_inst_ack_0, ack => convolution3D_CP_1120_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	150 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1271_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1271_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1271_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(156)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(156)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(156) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1271_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1271_inst_ack_1, ack => convolution3D_CP_1120_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	150 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1281_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1281_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1281_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(157)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(157)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(157) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1281_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1281_inst_ack_0, ack => convolution3D_CP_1120_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	150 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	161 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1281_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1281_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1281_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(158)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(158)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(158) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1281_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1281_inst_ack_1, ack => convolution3D_CP_1120_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	150 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1290_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1290_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1290_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(159)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(159)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(159) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1290_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1290_inst_ack_0, ack => convolution3D_CP_1120_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	150 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1290_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1290_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/type_cast_1290_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(160)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(160)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(160) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1290_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1290_inst_ack_1, ack => convolution3D_CP_1120_elements(160)); -- 
    -- CP-element group 161:  join  transition  place  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	154 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	158 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	244 
    -- CP-element group 161:  members (6) 
      -- CP-element group 161: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296/$exit
      -- CP-element group 161: 	 branch_block_stmt_435/assign_stmt_1238_to_assign_stmt_1296__exit__
      -- CP-element group 161: 	 branch_block_stmt_435/ifx_xend107_whilex_xbody
      -- CP-element group 161: 	 branch_block_stmt_435/ifx_xend107_whilex_xbody_PhiReq/$entry
      -- CP-element group 161: 	 branch_block_stmt_435/ifx_xend107_whilex_xbody_PhiReq/phi_stmt_1299/$entry
      -- CP-element group 161: 	 branch_block_stmt_435/ifx_xend107_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(161)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(161)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(161) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(152) & convolution3D_CP_1120_elements(154) & convolution3D_CP_1120_elements(156) & convolution3D_CP_1120_elements(158) & convolution3D_CP_1120_elements(160);
      gj_convolution3D_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	249 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1319_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1319_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1319_Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(162)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(162)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(162) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1319_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1319_inst_ack_0, ack => convolution3D_CP_1120_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	249 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	166 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1319_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1319_Update/ca
      -- CP-element group 163: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1319_Update/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(163)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(163)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(163) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1319_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1319_inst_ack_1, ack => convolution3D_CP_1120_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	249 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1323_Sample/ra
      -- CP-element group 164: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1323_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1323_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(164)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(164)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(164) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1323_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1323_inst_ack_0, ack => convolution3D_CP_1120_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	249 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1323_Update/ca
      -- CP-element group 165: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1323_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1323_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(165)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(165)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(165) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1323_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1323_inst_ack_1, ack => convolution3D_CP_1120_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	163 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1327_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1327_Sample/crr
      -- CP-element group 166: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1327_sample_start_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(166)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(166)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(166) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1327_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_2624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(166), ack => call_stmt_1327_call_req_0); -- 
    convolution3D_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(163) & convolution3D_CP_1120_elements(165);
      gj_convolution3D_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1327_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1327_Sample/cra
      -- CP-element group 167: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1327_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(167)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(167)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(167) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1327_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_2625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1327_call_ack_0, ack => convolution3D_CP_1120_elements(167)); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	249 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	171 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1327_Update/cca
      -- CP-element group 168: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1327_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1327_Update/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(168)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(168)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(168) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1327_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_2630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1327_call_ack_1, ack => convolution3D_CP_1120_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	249 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1334_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1334_Sample/cra
      -- CP-element group 169: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1334_Sample/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(169)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(169)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(169) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1334_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_2639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1334_call_ack_0, ack => convolution3D_CP_1120_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	249 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1334_Update/cca
      -- CP-element group 170: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1334_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1334_update_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(170)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(170)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(170) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1334_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_2644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1334_call_ack_1, ack => convolution3D_CP_1120_elements(170)); -- 
    -- CP-element group 171:  branch  join  transition  place  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	168 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (10) 
      -- CP-element group 171: 	 branch_block_stmt_435/R_exitcond7_1347_place
      -- CP-element group 171: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345__exit__
      -- CP-element group 171: 	 branch_block_stmt_435/if_stmt_1346__entry__
      -- CP-element group 171: 	 branch_block_stmt_435/if_stmt_1346_dead_link/$entry
      -- CP-element group 171: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/$exit
      -- CP-element group 171: 	 branch_block_stmt_435/if_stmt_1346_else_link/$entry
      -- CP-element group 171: 	 branch_block_stmt_435/if_stmt_1346_if_link/$entry
      -- CP-element group 171: 	 branch_block_stmt_435/if_stmt_1346_eval_test/branch_req
      -- CP-element group 171: 	 branch_block_stmt_435/if_stmt_1346_eval_test/$exit
      -- CP-element group 171: 	 branch_block_stmt_435/if_stmt_1346_eval_test/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(171)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(171)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(171) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_1346_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_2652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(171), ack => if_stmt_1346_branch_req_0); -- 
    convolution3D_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(168) & convolution3D_CP_1120_elements(170);
      gj_convolution3D_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: 	175 
    -- CP-element group 172:  members (18) 
      -- CP-element group 172: 	 branch_block_stmt_435/whilex_xbody_whilex_xend
      -- CP-element group 172: 	 branch_block_stmt_435/merge_stmt_1352__exit__
      -- CP-element group 172: 	 branch_block_stmt_435/assign_stmt_1357__entry__
      -- CP-element group 172: 	 branch_block_stmt_435/assign_stmt_1357/type_cast_1356_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_435/assign_stmt_1357/type_cast_1356_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_435/assign_stmt_1357/type_cast_1356_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_435/assign_stmt_1357/type_cast_1356_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_435/assign_stmt_1357/type_cast_1356_update_start_
      -- CP-element group 172: 	 branch_block_stmt_435/assign_stmt_1357/type_cast_1356_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_435/assign_stmt_1357/$entry
      -- CP-element group 172: 	 branch_block_stmt_435/if_stmt_1346_if_link/if_choice_transition
      -- CP-element group 172: 	 branch_block_stmt_435/if_stmt_1346_if_link/$exit
      -- CP-element group 172: 	 branch_block_stmt_435/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 172: 	 branch_block_stmt_435/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 172: 	 branch_block_stmt_435/merge_stmt_1352_PhiReqMerge
      -- CP-element group 172: 	 branch_block_stmt_435/merge_stmt_1352_PhiAck/$entry
      -- CP-element group 172: 	 branch_block_stmt_435/merge_stmt_1352_PhiAck/$exit
      -- CP-element group 172: 	 branch_block_stmt_435/merge_stmt_1352_PhiAck/dummy
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(172)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(172)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(172) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_1346_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1356_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1356_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_2657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1346_branch_ack_1, ack => convolution3D_CP_1120_elements(172)); -- 
    cr_2679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(172), ack => type_cast_1356_inst_req_1); -- 
    rr_2674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(172), ack => type_cast_1356_inst_req_0); -- 
    -- CP-element group 173:  fork  transition  place  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	245 
    -- CP-element group 173: 	246 
    -- CP-element group 173:  members (12) 
      -- CP-element group 173: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody
      -- CP-element group 173: 	 branch_block_stmt_435/if_stmt_1346_else_link/else_choice_transition
      -- CP-element group 173: 	 branch_block_stmt_435/if_stmt_1346_else_link/$exit
      -- CP-element group 173: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- CP-element group 173: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/$entry
      -- CP-element group 173: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/$entry
      -- CP-element group 173: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/type_cast_1302/$entry
      -- CP-element group 173: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/type_cast_1302/SplitProtocol/$entry
      -- CP-element group 173: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/type_cast_1302/SplitProtocol/Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/type_cast_1302/SplitProtocol/Sample/rr
      -- CP-element group 173: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/type_cast_1302/SplitProtocol/Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/type_cast_1302/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(173)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(173)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(173) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_1346_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1302_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1302_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_2661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1346_branch_ack_0, ack => convolution3D_CP_1120_elements(173)); -- 
    rr_3235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(173), ack => type_cast_1302_inst_req_0); -- 
    cr_3240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(173), ack => type_cast_1302_inst_req_1); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_435/assign_stmt_1357/type_cast_1356_Sample/ra
      -- CP-element group 174: 	 branch_block_stmt_435/assign_stmt_1357/type_cast_1356_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_435/assign_stmt_1357/type_cast_1356_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(174)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(174)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(174) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1356_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1356_inst_ack_0, ack => convolution3D_CP_1120_elements(174)); -- 
    -- CP-element group 175:  fork  transition  place  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	172 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175: 	177 
    -- CP-element group 175: 	179 
    -- CP-element group 175:  members (16) 
      -- CP-element group 175: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/call_stmt_1360_Update/ccr
      -- CP-element group 175: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/call_stmt_1360_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/type_cast_1364_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_435/assign_stmt_1357__exit__
      -- CP-element group 175: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373__entry__
      -- CP-element group 175: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/type_cast_1364_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/call_stmt_1360_Sample/crr
      -- CP-element group 175: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/call_stmt_1360_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/call_stmt_1360_update_start_
      -- CP-element group 175: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/call_stmt_1360_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/$entry
      -- CP-element group 175: 	 branch_block_stmt_435/assign_stmt_1357/type_cast_1356_Update/ca
      -- CP-element group 175: 	 branch_block_stmt_435/assign_stmt_1357/type_cast_1356_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_435/assign_stmt_1357/type_cast_1356_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_435/assign_stmt_1357/$exit
      -- CP-element group 175: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/type_cast_1364_update_start_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(175)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(175)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(175) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1356_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1360_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1364_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1360_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_2680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1356_inst_ack_1, ack => convolution3D_CP_1120_elements(175)); -- 
    ccr_2696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(175), ack => call_stmt_1360_call_req_1); -- 
    cr_2710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(175), ack => type_cast_1364_inst_req_1); -- 
    crr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(175), ack => call_stmt_1360_call_req_0); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/call_stmt_1360_Sample/cra
      -- CP-element group 176: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/call_stmt_1360_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/call_stmt_1360_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(176)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(176)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(176) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1360_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1360_call_ack_0, ack => convolution3D_CP_1120_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/call_stmt_1360_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/call_stmt_1360_Update/cca
      -- CP-element group 177: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/type_cast_1364_Sample/rr
      -- CP-element group 177: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/call_stmt_1360_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/type_cast_1364_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/type_cast_1364_sample_start_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(177)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(177)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(177) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1360_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1364_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_2697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1360_call_ack_1, ack => convolution3D_CP_1120_elements(177)); -- 
    rr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(177), ack => type_cast_1364_inst_req_0); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/type_cast_1364_Sample/ra
      -- CP-element group 178: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/type_cast_1364_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/type_cast_1364_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(178)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(178)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(178) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1364_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1364_inst_ack_0, ack => convolution3D_CP_1120_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	175 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/type_cast_1364_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/WPIPE_elapsed_time_pipe_1371_Sample/req
      -- CP-element group 179: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/WPIPE_elapsed_time_pipe_1371_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/WPIPE_elapsed_time_pipe_1371_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/type_cast_1364_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/type_cast_1364_Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(179)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(179)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(179) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1364_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:WPIPE_elapsed_time_pipe_1371_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_2711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1364_inst_ack_1, ack => convolution3D_CP_1120_elements(179)); -- 
    req_2719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(179), ack => WPIPE_elapsed_time_pipe_1371_inst_req_0); -- 
    -- CP-element group 180:  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/WPIPE_elapsed_time_pipe_1371_Update/req
      -- CP-element group 180: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/WPIPE_elapsed_time_pipe_1371_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/WPIPE_elapsed_time_pipe_1371_Sample/ack
      -- CP-element group 180: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/WPIPE_elapsed_time_pipe_1371_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/WPIPE_elapsed_time_pipe_1371_update_start_
      -- CP-element group 180: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/WPIPE_elapsed_time_pipe_1371_sample_completed_
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(180)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(180)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(180) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:WPIPE_elapsed_time_pipe_1371_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:WPIPE_elapsed_time_pipe_1371_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1371_inst_ack_0, ack => convolution3D_CP_1120_elements(180)); -- 
    req_2724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(180), ack => WPIPE_elapsed_time_pipe_1371_inst_req_1); -- 
    -- CP-element group 181:  transition  place  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (16) 
      -- CP-element group 181: 	 $exit
      -- CP-element group 181: 	 branch_block_stmt_435/$exit
      -- CP-element group 181: 	 branch_block_stmt_435/branch_block_stmt_435__exit__
      -- CP-element group 181: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373__exit__
      -- CP-element group 181: 	 branch_block_stmt_435/return__
      -- CP-element group 181: 	 branch_block_stmt_435/merge_stmt_1376__exit__
      -- CP-element group 181: 	 branch_block_stmt_435/merge_stmt_1376_PhiReqMerge
      -- CP-element group 181: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/WPIPE_elapsed_time_pipe_1371_Update/ack
      -- CP-element group 181: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/$exit
      -- CP-element group 181: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/WPIPE_elapsed_time_pipe_1371_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_435/call_stmt_1360_to_assign_stmt_1373/WPIPE_elapsed_time_pipe_1371_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_435/return___PhiReq/$entry
      -- CP-element group 181: 	 branch_block_stmt_435/return___PhiReq/$exit
      -- CP-element group 181: 	 branch_block_stmt_435/merge_stmt_1376_PhiAck/$entry
      -- CP-element group 181: 	 branch_block_stmt_435/merge_stmt_1376_PhiAck/$exit
      -- CP-element group 181: 	 branch_block_stmt_435/merge_stmt_1376_PhiAck/dummy
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(181)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(181)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(181) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:WPIPE_elapsed_time_pipe_1371_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1371_inst_ack_1, ack => convolution3D_CP_1120_elements(181)); -- 
    -- CP-element group 182:  transition  output  delay-element  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	36 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	186 
    -- CP-element group 182:  members (5) 
      -- CP-element group 182: 	 branch_block_stmt_435/bbx_xnph197_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_req
      -- CP-element group 182: 	 branch_block_stmt_435/bbx_xnph197_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/type_cast_579_konst_delay_trans
      -- CP-element group 182: 	 branch_block_stmt_435/bbx_xnph197_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/$exit
      -- CP-element group 182: 	 branch_block_stmt_435/bbx_xnph197_forx_xbody_PhiReq/phi_stmt_575/$exit
      -- CP-element group 182: 	 branch_block_stmt_435/bbx_xnph197_forx_xbody_PhiReq/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(182)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(182)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(182) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_575_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_575_req_2748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_575_req_2748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(182), ack => phi_stmt_575_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(182) is a control-delay.
    cp_element_182_delay: control_delay_element  generic map(name => " 182_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(36), ack => convolution3D_CP_1120_elements(182), clk => clk, reset =>reset);
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	62 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/type_cast_581/SplitProtocol/Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/type_cast_581/SplitProtocol/Sample/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(183)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(183)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(183) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_581_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_581_inst_ack_0, ack => convolution3D_CP_1120_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	62 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (2) 
      -- CP-element group 184: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/type_cast_581/SplitProtocol/Update/ca
      -- CP-element group 184: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/type_cast_581/SplitProtocol/Update/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(184)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(184)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(184) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_581_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_581_inst_ack_1, ack => convolution3D_CP_1120_elements(184)); -- 
    -- CP-element group 185:  join  transition  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 185: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_req
      -- CP-element group 185: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/$exit
      -- CP-element group 185: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/type_cast_581/SplitProtocol/$exit
      -- CP-element group 185: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/$exit
      -- CP-element group 185: 	 branch_block_stmt_435/forx_xbody_forx_xbody_PhiReq/phi_stmt_575/phi_stmt_575_sources/type_cast_581/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(185)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(185)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(185) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_575_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_575_req_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_575_req_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(185), ack => phi_stmt_575_req_1); -- 
    convolution3D_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(183) & convolution3D_CP_1120_elements(184);
      gj_convolution3D_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  merge  transition  place  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	182 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (2) 
      -- CP-element group 186: 	 branch_block_stmt_435/merge_stmt_574_PhiReqMerge
      -- CP-element group 186: 	 branch_block_stmt_435/merge_stmt_574_PhiAck/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(186)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(186)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(186) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_CP_1120_elements(186) <= OrReduce(convolution3D_CP_1120_elements(182) & convolution3D_CP_1120_elements(185));
    -- CP-element group 187:  fork  transition  place  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	37 
    -- CP-element group 187: 	38 
    -- CP-element group 187: 	40 
    -- CP-element group 187: 	41 
    -- CP-element group 187: 	44 
    -- CP-element group 187: 	48 
    -- CP-element group 187: 	52 
    -- CP-element group 187: 	56 
    -- CP-element group 187: 	59 
    -- CP-element group 187:  members (44) 
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Update/word_access_complete/word_0/cr
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_index_scale_1/$exit
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_608_Update/cr
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_591_Sample/rr
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_608_update_start_
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Update/word_access_complete/word_0/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_index_scale_1/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_index_resize_1/index_resize_ack
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_626_update_start_
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_index_resize_1/index_resize_req
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Update/word_access_complete/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_index_resize_1/$exit
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_index_resize_1/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/addr_of_588_complete/req
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_608_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_index_computed_1
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/addr_of_588_complete/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_index_resized_1
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_591_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_595_update_start_
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_index_scale_1/scale_rename_req
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/addr_of_588_update_start_
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_595_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_595_Update/cr
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_index_scale_1/scale_rename_ack
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_index_scaled_1
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_644_Update/cr
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_644_update_start_
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_final_index_sum_regn_update_start
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_final_index_sum_regn_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_final_index_sum_regn_Sample/req
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_final_index_sum_regn_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/array_obj_ref_587_final_index_sum_regn_Update/req
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_626_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/RPIPE_maxpool_input_pipe_591_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/merge_stmt_574_PhiAck/phi_stmt_575_ack
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/ptr_deref_652_update_start_
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_626_Update/cr
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665/type_cast_644_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_435/merge_stmt_574__exit__
      -- CP-element group 187: 	 branch_block_stmt_435/assign_stmt_589_to_assign_stmt_665__entry__
      -- CP-element group 187: 	 branch_block_stmt_435/merge_stmt_574_PhiAck/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(187)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(187)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(187) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_575_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_652_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_608_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_591_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_588_final_reg_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_595_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_644_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_587_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_587_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_626_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_575_ack_2779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_575_ack_0, ack => convolution3D_CP_1120_elements(187)); -- 
    cr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(187), ack => ptr_deref_652_store_0_req_1); -- 
    cr_1578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(187), ack => type_cast_608_inst_req_1); -- 
    rr_1531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(187), ack => RPIPE_maxpool_input_pipe_591_inst_req_0); -- 
    req_1522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(187), ack => addr_of_588_final_reg_req_1); -- 
    cr_1550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(187), ack => type_cast_595_inst_req_1); -- 
    cr_1634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(187), ack => type_cast_644_inst_req_1); -- 
    req_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(187), ack => array_obj_ref_587_index_offset_req_0); -- 
    req_1507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(187), ack => array_obj_ref_587_index_offset_req_1); -- 
    cr_1606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(187), ack => type_cast_626_inst_req_1); -- 
    -- CP-element group 188:  transition  output  delay-element  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	25 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	192 
    -- CP-element group 188:  members (5) 
      -- CP-element group 188: 	 branch_block_stmt_435/entry_forx_xend_PhiReq/$exit
      -- CP-element group 188: 	 branch_block_stmt_435/entry_forx_xend_PhiReq/phi_stmt_697/$exit
      -- CP-element group 188: 	 branch_block_stmt_435/entry_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/$exit
      -- CP-element group 188: 	 branch_block_stmt_435/entry_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/type_cast_703_konst_delay_trans
      -- CP-element group 188: 	 branch_block_stmt_435/entry_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(188)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(188)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(188) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_697_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_697_req_2802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_697_req_2802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(188), ack => phi_stmt_697_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(188) is a control-delay.
    cp_element_188_delay: control_delay_element  generic map(name => " 188_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(25), ack => convolution3D_CP_1120_elements(188), clk => clk, reset =>reset);
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	61 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (2) 
      -- CP-element group 189: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/type_cast_700/SplitProtocol/Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/type_cast_700/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(189)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(189)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(189) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_700_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_700_inst_ack_0, ack => convolution3D_CP_1120_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	61 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (2) 
      -- CP-element group 190: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/type_cast_700/SplitProtocol/Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/type_cast_700/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(190)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(190)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(190) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_700_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_700_inst_ack_1, ack => convolution3D_CP_1120_elements(190)); -- 
    -- CP-element group 191:  join  transition  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 191: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/$exit
      -- CP-element group 191: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/$exit
      -- CP-element group 191: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/type_cast_700/$exit
      -- CP-element group 191: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_sources/type_cast_700/SplitProtocol/$exit
      -- CP-element group 191: 	 branch_block_stmt_435/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_697/phi_stmt_697_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(191)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(191)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(191) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_697_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_697_req_2828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_697_req_2828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(191), ack => phi_stmt_697_req_0); -- 
    convolution3D_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(189) & convolution3D_CP_1120_elements(190);
      gj_convolution3D_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  merge  transition  place  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	188 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (2) 
      -- CP-element group 192: 	 branch_block_stmt_435/merge_stmt_696_PhiReqMerge
      -- CP-element group 192: 	 branch_block_stmt_435/merge_stmt_696_PhiAck/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(192)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(192)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(192) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_CP_1120_elements(192) <= OrReduce(convolution3D_CP_1120_elements(188) & convolution3D_CP_1120_elements(191));
    -- CP-element group 193:  branch  transition  place  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	63 
    -- CP-element group 193: 	64 
    -- CP-element group 193:  members (15) 
      -- CP-element group 193: 	 branch_block_stmt_435/R_tobool_718_place
      -- CP-element group 193: 	 branch_block_stmt_435/assign_stmt_710_to_assign_stmt_716/$entry
      -- CP-element group 193: 	 branch_block_stmt_435/if_stmt_717_eval_test/$entry
      -- CP-element group 193: 	 branch_block_stmt_435/if_stmt_717_if_link/$entry
      -- CP-element group 193: 	 branch_block_stmt_435/if_stmt_717_eval_test/$exit
      -- CP-element group 193: 	 branch_block_stmt_435/if_stmt_717_eval_test/branch_req
      -- CP-element group 193: 	 branch_block_stmt_435/if_stmt_717_else_link/$entry
      -- CP-element group 193: 	 branch_block_stmt_435/if_stmt_717_dead_link/$entry
      -- CP-element group 193: 	 branch_block_stmt_435/assign_stmt_710_to_assign_stmt_716/$exit
      -- CP-element group 193: 	 branch_block_stmt_435/merge_stmt_696__exit__
      -- CP-element group 193: 	 branch_block_stmt_435/assign_stmt_710_to_assign_stmt_716__entry__
      -- CP-element group 193: 	 branch_block_stmt_435/assign_stmt_710_to_assign_stmt_716__exit__
      -- CP-element group 193: 	 branch_block_stmt_435/if_stmt_717__entry__
      -- CP-element group 193: 	 branch_block_stmt_435/merge_stmt_696_PhiAck/$exit
      -- CP-element group 193: 	 branch_block_stmt_435/merge_stmt_696_PhiAck/phi_stmt_697_ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(193)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(193)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(193) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_697_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_717_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_697_ack_2833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_697_ack_0, ack => convolution3D_CP_1120_elements(193)); -- 
    branch_req_1718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(193), ack => if_stmt_717_branch_req_0); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	74 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (2) 
      -- CP-element group 194: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_747/SplitProtocol/Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_747/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(194)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(194)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(194) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_747_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_747_inst_ack_0, ack => convolution3D_CP_1120_elements(194)); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	74 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (2) 
      -- CP-element group 195: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_747/SplitProtocol/Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_747/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(195)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(195)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(195) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_747_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_747_inst_ack_1, ack => convolution3D_CP_1120_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	200 
    -- CP-element group 196:  members (5) 
      -- CP-element group 196: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/$exit
      -- CP-element group 196: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/$exit
      -- CP-element group 196: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_747/$exit
      -- CP-element group 196: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_747/SplitProtocol/$exit
      -- CP-element group 196: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(196)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(196)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(196) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_744_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_744_req_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_744_req_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(196), ack => phi_stmt_744_req_0); -- 
    convolution3D_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(194) & convolution3D_CP_1120_elements(195);
      gj_convolution3D_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	74 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (2) 
      -- CP-element group 197: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(197)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(197)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(197) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_754_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_754_inst_ack_0, ack => convolution3D_CP_1120_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	74 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (2) 
      -- CP-element group 198: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(198)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(198)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(198) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_754_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_754_inst_ack_1, ack => convolution3D_CP_1120_elements(198)); -- 
    -- CP-element group 199:  join  transition  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (5) 
      -- CP-element group 199: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/$exit
      -- CP-element group 199: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/$exit
      -- CP-element group 199: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/$exit
      -- CP-element group 199: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/$exit
      -- CP-element group 199: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(199)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(199)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(199) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_751_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_751_req_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_751_req_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(199), ack => phi_stmt_751_req_0); -- 
    convolution3D_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(197) & convolution3D_CP_1120_elements(198);
      gj_convolution3D_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  join  transition  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	196 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	204 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_435/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(200)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(200)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(200) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(196) & convolution3D_CP_1120_elements(199);
      gj_convolution3D_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  transition  output  delay-element  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	68 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	203 
    -- CP-element group 201:  members (4) 
      -- CP-element group 201: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_744/$exit
      -- CP-element group 201: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/$exit
      -- CP-element group 201: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_750_konst_delay_trans
      -- CP-element group 201: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_744/phi_stmt_744_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(201)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(201)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(201) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_744_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_744_req_2905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_744_req_2905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(201), ack => phi_stmt_744_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(201) is a control-delay.
    cp_element_201_delay: control_delay_element  generic map(name => " 201_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(68), ack => convolution3D_CP_1120_elements(201), clk => clk, reset =>reset);
    -- CP-element group 202:  transition  output  delay-element  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	68 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (4) 
      -- CP-element group 202: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_751/$exit
      -- CP-element group 202: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/$exit
      -- CP-element group 202: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_757_konst_delay_trans
      -- CP-element group 202: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_751/phi_stmt_751_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(202)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(202)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(202) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_751_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_751_req_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_751_req_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(202), ack => phi_stmt_751_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(202) is a control-delay.
    cp_element_202_delay: control_delay_element  generic map(name => " 202_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(68), ack => convolution3D_CP_1120_elements(202), clk => clk, reset =>reset);
    -- CP-element group 203:  join  transition  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	201 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_435/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(203)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(203)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(203) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(201) & convolution3D_CP_1120_elements(202);
      gj_convolution3D_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  merge  fork  transition  place  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	200 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (2) 
      -- CP-element group 204: 	 branch_block_stmt_435/merge_stmt_743_PhiReqMerge
      -- CP-element group 204: 	 branch_block_stmt_435/merge_stmt_743_PhiAck/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(204)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(204)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(204) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_CP_1120_elements(204) <= OrReduce(convolution3D_CP_1120_elements(200) & convolution3D_CP_1120_elements(203));
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	207 
    -- CP-element group 205:  members (1) 
      -- CP-element group 205: 	 branch_block_stmt_435/merge_stmt_743_PhiAck/phi_stmt_744_ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(205)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(205)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(205) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_744_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_744_ack_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_744_ack_0, ack => convolution3D_CP_1120_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 branch_block_stmt_435/merge_stmt_743_PhiAck/phi_stmt_751_ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(206)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(206)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(206) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_751_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_751_ack_2919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_751_ack_0, ack => convolution3D_CP_1120_elements(206)); -- 
    -- CP-element group 207:  join  fork  transition  place  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	205 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	69 
    -- CP-element group 207: 	72 
    -- CP-element group 207:  members (10) 
      -- CP-element group 207: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/RPIPE_maxpool_input_pipe_760_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/$entry
      -- CP-element group 207: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/type_cast_764_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/type_cast_764_Update/cr
      -- CP-element group 207: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/type_cast_764_update_start_
      -- CP-element group 207: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/RPIPE_maxpool_input_pipe_760_Sample/rr
      -- CP-element group 207: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787/RPIPE_maxpool_input_pipe_760_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_435/merge_stmt_743__exit__
      -- CP-element group 207: 	 branch_block_stmt_435/assign_stmt_761_to_assign_stmt_787__entry__
      -- CP-element group 207: 	 branch_block_stmt_435/merge_stmt_743_PhiAck/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(207)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(207)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(207) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_764_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_760_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cr_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(207), ack => type_cast_764_inst_req_1); -- 
    rr_1771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(207), ack => RPIPE_maxpool_input_pipe_760_inst_req_0); -- 
    convolution3D_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(205) & convolution3D_CP_1120_elements(206);
      gj_convolution3D_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	73 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (2) 
      -- CP-element group 208: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/type_cast_798/SplitProtocol/Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/type_cast_798/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(208)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(208)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(208) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_798_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_798_inst_ack_0, ack => convolution3D_CP_1120_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	73 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (2) 
      -- CP-element group 209: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/type_cast_798/SplitProtocol/Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/type_cast_798/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(209)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(209)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(209) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_798_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_798_inst_ack_1, ack => convolution3D_CP_1120_elements(209)); -- 
    -- CP-element group 210:  join  transition  place  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (8) 
      -- CP-element group 210: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- CP-element group 210: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/$exit
      -- CP-element group 210: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/$exit
      -- CP-element group 210: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/type_cast_798/$exit
      -- CP-element group 210: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_sources/type_cast_798/SplitProtocol/$exit
      -- CP-element group 210: 	 branch_block_stmt_435/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_795/phi_stmt_795_req
      -- CP-element group 210: 	 branch_block_stmt_435/merge_stmt_794_PhiReqMerge
      -- CP-element group 210: 	 branch_block_stmt_435/merge_stmt_794_PhiAck/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(210)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(210)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(210) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_795_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_795_req_2949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_795_req_2949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(210), ack => phi_stmt_795_req_0); -- 
    convolution3D_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(208) & convolution3D_CP_1120_elements(209);
      gj_convolution3D_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	75 
    -- CP-element group 211: 	76 
    -- CP-element group 211: 	78 
    -- CP-element group 211: 	80 
    -- CP-element group 211:  members (29) 
      -- CP-element group 211: 	 branch_block_stmt_435/merge_stmt_794__exit__
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833__entry__
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/$entry
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/addr_of_828_update_start_
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_index_resized_1
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_index_scaled_1
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_index_computed_1
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_index_resize_1/$entry
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_index_resize_1/$exit
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_index_resize_1/index_resize_req
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_index_resize_1/index_resize_ack
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_index_scale_1/$entry
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_index_scale_1/$exit
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_index_scale_1/scale_rename_req
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_index_scale_1/scale_rename_ack
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_final_index_sum_regn_update_start
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_final_index_sum_regn_Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_final_index_sum_regn_Sample/req
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_final_index_sum_regn_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/array_obj_ref_827_final_index_sum_regn_Update/req
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/addr_of_828_complete/$entry
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/addr_of_828_complete/req
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_update_start_
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Update/word_access_complete/$entry
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Update/word_access_complete/word_0/$entry
      -- CP-element group 211: 	 branch_block_stmt_435/assign_stmt_805_to_assign_stmt_833/ptr_deref_831_Update/word_access_complete/word_0/cr
      -- CP-element group 211: 	 branch_block_stmt_435/merge_stmt_794_PhiAck/$exit
      -- CP-element group 211: 	 branch_block_stmt_435/merge_stmt_794_PhiAck/phi_stmt_795_ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(211)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(211)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(211) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_795_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_827_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_827_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_828_final_reg_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_831_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_795_ack_2954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_795_ack_0, ack => convolution3D_CP_1120_elements(211)); -- 
    req_1838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(211), ack => array_obj_ref_827_index_offset_req_0); -- 
    req_1843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(211), ack => array_obj_ref_827_index_offset_req_1); -- 
    req_1858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(211), ack => addr_of_828_final_reg_req_1); -- 
    cr_1908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(211), ack => ptr_deref_831_store_0_req_1); -- 
    -- CP-element group 212:  merge  fork  transition  place  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	63 
    -- CP-element group 212: 	81 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	82 
    -- CP-element group 212: 	83 
    -- CP-element group 212: 	84 
    -- CP-element group 212: 	85 
    -- CP-element group 212: 	86 
    -- CP-element group 212: 	87 
    -- CP-element group 212:  members (25) 
      -- CP-element group 212: 	 branch_block_stmt_435/merge_stmt_835__exit__
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883__entry__
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/$entry
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_838_sample_start_
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_838_update_start_
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_838_Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_838_Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_838_Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_838_Update/cr
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_842_sample_start_
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_842_update_start_
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_842_Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_842_Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_842_Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_842_Update/cr
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_846_sample_start_
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_846_update_start_
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_846_Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_846_Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_846_Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_435/assign_stmt_839_to_assign_stmt_883/type_cast_846_Update/cr
      -- CP-element group 212: 	 branch_block_stmt_435/merge_stmt_835_PhiReqMerge
      -- CP-element group 212: 	 branch_block_stmt_435/merge_stmt_835_PhiAck/$entry
      -- CP-element group 212: 	 branch_block_stmt_435/merge_stmt_835_PhiAck/$exit
      -- CP-element group 212: 	 branch_block_stmt_435/merge_stmt_835_PhiAck/dummy
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(212)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(212)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(212) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_838_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_838_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_842_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_842_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_846_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_846_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    rr_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(212), ack => type_cast_838_inst_req_0); -- 
    cr_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(212), ack => type_cast_838_inst_req_1); -- 
    rr_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(212), ack => type_cast_842_inst_req_0); -- 
    cr_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(212), ack => type_cast_842_inst_req_1); -- 
    rr_1948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(212), ack => type_cast_846_inst_req_0); -- 
    cr_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(212), ack => type_cast_846_inst_req_1); -- 
    convolution3D_CP_1120_elements(212) <= OrReduce(convolution3D_CP_1120_elements(63) & convolution3D_CP_1120_elements(81));
    -- CP-element group 213:  transition  output  delay-element  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	103 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	217 
    -- CP-element group 213:  members (5) 
      -- CP-element group 213: 	 branch_block_stmt_435/bbx_xnph_forx_xbody67_PhiReq/$exit
      -- CP-element group 213: 	 branch_block_stmt_435/bbx_xnph_forx_xbody67_PhiReq/phi_stmt_964/$exit
      -- CP-element group 213: 	 branch_block_stmt_435/bbx_xnph_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/$exit
      -- CP-element group 213: 	 branch_block_stmt_435/bbx_xnph_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/type_cast_968_konst_delay_trans
      -- CP-element group 213: 	 branch_block_stmt_435/bbx_xnph_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(213)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(213)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(213) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_964_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_964_req_2988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_964_req_2988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(213), ack => phi_stmt_964_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(213) is a control-delay.
    cp_element_213_delay: control_delay_element  generic map(name => " 213_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(103), ack => convolution3D_CP_1120_elements(213), clk => clk, reset =>reset);
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	129 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (2) 
      -- CP-element group 214: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/type_cast_970/SplitProtocol/Sample/$exit
      -- CP-element group 214: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/type_cast_970/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(214)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(214)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(214) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_970_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_970_inst_ack_0, ack => convolution3D_CP_1120_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	129 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (2) 
      -- CP-element group 215: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/type_cast_970/SplitProtocol/Update/$exit
      -- CP-element group 215: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/type_cast_970/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(215)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(215)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(215) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_970_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_970_inst_ack_1, ack => convolution3D_CP_1120_elements(215)); -- 
    -- CP-element group 216:  join  transition  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (6) 
      -- CP-element group 216: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/$exit
      -- CP-element group 216: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/$exit
      -- CP-element group 216: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/$exit
      -- CP-element group 216: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/type_cast_970/$exit
      -- CP-element group 216: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_sources/type_cast_970/SplitProtocol/$exit
      -- CP-element group 216: 	 branch_block_stmt_435/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_964/phi_stmt_964_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(216)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(216)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(216) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_964_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_964_req_3014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_964_req_3014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(216), ack => phi_stmt_964_req_1); -- 
    convolution3D_cp_element_group_216: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_216"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(214) & convolution3D_CP_1120_elements(215);
      gj_convolution3D_cp_element_group_216 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 217:  merge  transition  place  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	213 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (2) 
      -- CP-element group 217: 	 branch_block_stmt_435/merge_stmt_963_PhiReqMerge
      -- CP-element group 217: 	 branch_block_stmt_435/merge_stmt_963_PhiAck/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(217)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(217)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(217) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_CP_1120_elements(217) <= OrReduce(convolution3D_CP_1120_elements(213) & convolution3D_CP_1120_elements(216));
    -- CP-element group 218:  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	104 
    -- CP-element group 218: 	105 
    -- CP-element group 218: 	107 
    -- CP-element group 218: 	108 
    -- CP-element group 218: 	111 
    -- CP-element group 218: 	115 
    -- CP-element group 218: 	119 
    -- CP-element group 218: 	123 
    -- CP-element group 218: 	126 
    -- CP-element group 218:  members (44) 
      -- CP-element group 218: 	 branch_block_stmt_435/merge_stmt_963__exit__
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054__entry__
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/addr_of_977_update_start_
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_index_resized_1
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_index_scaled_1
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_index_computed_1
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_index_resize_1/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_index_resize_1/$exit
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_index_resize_1/index_resize_req
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_index_resize_1/index_resize_ack
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_index_scale_1/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_index_scale_1/$exit
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_index_scale_1/scale_rename_req
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_index_scale_1/scale_rename_ack
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_final_index_sum_regn_update_start
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_final_index_sum_regn_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_final_index_sum_regn_Sample/req
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_final_index_sum_regn_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/array_obj_ref_976_final_index_sum_regn_Update/req
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/addr_of_977_complete/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/addr_of_977_complete/req
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_980_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_980_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/RPIPE_maxpool_input_pipe_980_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_984_update_start_
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_984_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_984_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_997_update_start_
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_997_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_997_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1015_update_start_
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1015_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1015_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1033_update_start_
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1033_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/type_cast_1033_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_update_start_
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Update/word_access_complete/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Update/word_access_complete/word_0/$entry
      -- CP-element group 218: 	 branch_block_stmt_435/assign_stmt_978_to_assign_stmt_1054/ptr_deref_1041_Update/word_access_complete/word_0/cr
      -- CP-element group 218: 	 branch_block_stmt_435/merge_stmt_963_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_435/merge_stmt_963_PhiAck/phi_stmt_964_ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(218)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(218)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(218) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_964_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_976_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_976_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_977_final_reg_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_980_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_984_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_997_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1015_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1033_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_1041_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_964_ack_3019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_964_ack_0, ack => convolution3D_CP_1120_elements(218)); -- 
    req_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(218), ack => array_obj_ref_976_index_offset_req_0); -- 
    req_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(218), ack => array_obj_ref_976_index_offset_req_1); -- 
    req_2108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(218), ack => addr_of_977_final_reg_req_1); -- 
    rr_2117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(218), ack => RPIPE_maxpool_input_pipe_980_inst_req_0); -- 
    cr_2136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(218), ack => type_cast_984_inst_req_1); -- 
    cr_2164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(218), ack => type_cast_997_inst_req_1); -- 
    cr_2192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(218), ack => type_cast_1015_inst_req_1); -- 
    cr_2220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(218), ack => type_cast_1033_inst_req_1); -- 
    cr_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(218), ack => ptr_deref_1041_store_0_req_1); -- 
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	128 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (2) 
      -- CP-element group 219: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/type_cast_1089/SplitProtocol/Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/type_cast_1089/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(219)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(219)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(219) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1089_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1089_inst_ack_0, ack => convolution3D_CP_1120_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	128 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220:  members (2) 
      -- CP-element group 220: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/type_cast_1089/SplitProtocol/Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/type_cast_1089/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(220)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(220)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(220) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1089_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1089_inst_ack_1, ack => convolution3D_CP_1120_elements(220)); -- 
    -- CP-element group 221:  join  transition  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (6) 
      -- CP-element group 221: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/$exit
      -- CP-element group 221: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/$exit
      -- CP-element group 221: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/$exit
      -- CP-element group 221: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/type_cast_1089/$exit
      -- CP-element group 221: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/type_cast_1089/SplitProtocol/$exit
      -- CP-element group 221: 	 branch_block_stmt_435/forx_xcond60x_xforx_xend95_crit_edge_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(221)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(221)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(221) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1086_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1086_req_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1086_req_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(221), ack => phi_stmt_1086_req_0); -- 
    convolution3D_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(219) & convolution3D_CP_1120_elements(220);
      gj_convolution3D_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  transition  output  delay-element  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	90 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (5) 
      -- CP-element group 222: 	 branch_block_stmt_435/ifx_xend_forx_xend95_PhiReq/$exit
      -- CP-element group 222: 	 branch_block_stmt_435/ifx_xend_forx_xend95_PhiReq/phi_stmt_1086/$exit
      -- CP-element group 222: 	 branch_block_stmt_435/ifx_xend_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/$exit
      -- CP-element group 222: 	 branch_block_stmt_435/ifx_xend_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_sources/type_cast_1092_konst_delay_trans
      -- CP-element group 222: 	 branch_block_stmt_435/ifx_xend_forx_xend95_PhiReq/phi_stmt_1086/phi_stmt_1086_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(222)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(222)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(222) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1086_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1086_req_3068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1086_req_3068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(222), ack => phi_stmt_1086_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(222) is a control-delay.
    cp_element_222_delay: control_delay_element  generic map(name => " 222_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(90), ack => convolution3D_CP_1120_elements(222), clk => clk, reset =>reset);
    -- CP-element group 223:  merge  transition  place  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (2) 
      -- CP-element group 223: 	 branch_block_stmt_435/merge_stmt_1085_PhiReqMerge
      -- CP-element group 223: 	 branch_block_stmt_435/merge_stmt_1085_PhiAck/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(223)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(223)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(223) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_CP_1120_elements(223) <= OrReduce(convolution3D_CP_1120_elements(221) & convolution3D_CP_1120_elements(222));
    -- CP-element group 224:  branch  transition  place  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	130 
    -- CP-element group 224: 	131 
    -- CP-element group 224:  members (15) 
      -- CP-element group 224: 	 branch_block_stmt_435/if_stmt_1106_else_link/$entry
      -- CP-element group 224: 	 branch_block_stmt_435/merge_stmt_1085__exit__
      -- CP-element group 224: 	 branch_block_stmt_435/assign_stmt_1099_to_assign_stmt_1105__entry__
      -- CP-element group 224: 	 branch_block_stmt_435/assign_stmt_1099_to_assign_stmt_1105__exit__
      -- CP-element group 224: 	 branch_block_stmt_435/if_stmt_1106__entry__
      -- CP-element group 224: 	 branch_block_stmt_435/if_stmt_1106_if_link/$entry
      -- CP-element group 224: 	 branch_block_stmt_435/if_stmt_1106_eval_test/branch_req
      -- CP-element group 224: 	 branch_block_stmt_435/if_stmt_1106_eval_test/$exit
      -- CP-element group 224: 	 branch_block_stmt_435/if_stmt_1106_eval_test/$entry
      -- CP-element group 224: 	 branch_block_stmt_435/if_stmt_1106_dead_link/$entry
      -- CP-element group 224: 	 branch_block_stmt_435/assign_stmt_1099_to_assign_stmt_1105/$exit
      -- CP-element group 224: 	 branch_block_stmt_435/assign_stmt_1099_to_assign_stmt_1105/$entry
      -- CP-element group 224: 	 branch_block_stmt_435/R_tobool98_1107_place
      -- CP-element group 224: 	 branch_block_stmt_435/merge_stmt_1085_PhiAck/$exit
      -- CP-element group 224: 	 branch_block_stmt_435/merge_stmt_1085_PhiAck/phi_stmt_1086_ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(224)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(224)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(224) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1086_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:if_stmt_1106_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1086_ack_3073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1086_ack_0, ack => convolution3D_CP_1120_elements(224)); -- 
    branch_req_2304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(224), ack => if_stmt_1106_branch_req_0); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	141 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (2) 
      -- CP-element group 225: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/type_cast_1141/SplitProtocol/Sample/$exit
      -- CP-element group 225: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/type_cast_1141/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(225)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(225)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(225) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1141_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1141_inst_ack_0, ack => convolution3D_CP_1120_elements(225)); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	141 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (2) 
      -- CP-element group 226: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/type_cast_1141/SplitProtocol/Update/$exit
      -- CP-element group 226: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/type_cast_1141/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(226)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(226)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(226) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1141_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1141_inst_ack_1, ack => convolution3D_CP_1120_elements(226)); -- 
    -- CP-element group 227:  join  transition  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	231 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/$exit
      -- CP-element group 227: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/$exit
      -- CP-element group 227: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/type_cast_1141/$exit
      -- CP-element group 227: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/type_cast_1141/SplitProtocol/$exit
      -- CP-element group 227: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(227)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(227)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(227) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1138_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1138_req_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1138_req_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(227), ack => phi_stmt_1138_req_0); -- 
    convolution3D_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(225) & convolution3D_CP_1120_elements(226);
      gj_convolution3D_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	141 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (2) 
      -- CP-element group 228: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/type_cast_1148/SplitProtocol/Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/type_cast_1148/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(228)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(228)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(228) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1148_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1148_inst_ack_0, ack => convolution3D_CP_1120_elements(228)); -- 
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	141 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (2) 
      -- CP-element group 229: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/type_cast_1148/SplitProtocol/Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/type_cast_1148/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(229)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(229)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(229) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1148_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1148_inst_ack_1, ack => convolution3D_CP_1120_elements(229)); -- 
    -- CP-element group 230:  join  transition  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (5) 
      -- CP-element group 230: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/$exit
      -- CP-element group 230: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/$exit
      -- CP-element group 230: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/type_cast_1148/$exit
      -- CP-element group 230: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/type_cast_1148/SplitProtocol/$exit
      -- CP-element group 230: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(230)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(230)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(230) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1145_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1145_req_3134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1145_req_3134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(230), ack => phi_stmt_1145_req_0); -- 
    convolution3D_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(228) & convolution3D_CP_1120_elements(229);
      gj_convolution3D_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  join  transition  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	227 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	235 
    -- CP-element group 231:  members (1) 
      -- CP-element group 231: 	 branch_block_stmt_435/forx_xbodyx_xi181_forx_xbodyx_xi181_PhiReq/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(231)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(231)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(231) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(227) & convolution3D_CP_1120_elements(230);
      gj_convolution3D_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  transition  output  delay-element  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	135 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	234 
    -- CP-element group 232:  members (4) 
      -- CP-element group 232: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/$exit
      -- CP-element group 232: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/$exit
      -- CP-element group 232: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_sources/type_cast_1144_konst_delay_trans
      -- CP-element group 232: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/phi_stmt_1138/phi_stmt_1138_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(232)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(232)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(232) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1138_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1138_req_3145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1138_req_3145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(232), ack => phi_stmt_1138_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(232) is a control-delay.
    cp_element_232_delay: control_delay_element  generic map(name => " 232_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(135), ack => convolution3D_CP_1120_elements(232), clk => clk, reset =>reset);
    -- CP-element group 233:  transition  output  delay-element  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	135 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (4) 
      -- CP-element group 233: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/$exit
      -- CP-element group 233: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/$exit
      -- CP-element group 233: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_sources/type_cast_1151_konst_delay_trans
      -- CP-element group 233: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/phi_stmt_1145/phi_stmt_1145_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(233)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(233)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(233) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1145_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1145_req_3153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1145_req_3153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(233), ack => phi_stmt_1145_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(233) is a control-delay.
    cp_element_233_delay: control_delay_element  generic map(name => " 233_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(135), ack => convolution3D_CP_1120_elements(233), clk => clk, reset =>reset);
    -- CP-element group 234:  join  transition  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	232 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (1) 
      -- CP-element group 234: 	 branch_block_stmt_435/forx_xbodyx_xi181x_xpreheader_forx_xbodyx_xi181_PhiReq/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(234)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(234)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(234) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(232) & convolution3D_CP_1120_elements(233);
      gj_convolution3D_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  merge  fork  transition  place  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	231 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235: 	237 
    -- CP-element group 235:  members (2) 
      -- CP-element group 235: 	 branch_block_stmt_435/merge_stmt_1137_PhiReqMerge
      -- CP-element group 235: 	 branch_block_stmt_435/merge_stmt_1137_PhiAck/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(235)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(235)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(235) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_CP_1120_elements(235) <= OrReduce(convolution3D_CP_1120_elements(231) & convolution3D_CP_1120_elements(234));
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	238 
    -- CP-element group 236:  members (1) 
      -- CP-element group 236: 	 branch_block_stmt_435/merge_stmt_1137_PhiAck/phi_stmt_1138_ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(236)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(236)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(236) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1138_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1138_ack_3158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1138_ack_0, ack => convolution3D_CP_1120_elements(236)); -- 
    -- CP-element group 237:  transition  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	235 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (1) 
      -- CP-element group 237: 	 branch_block_stmt_435/merge_stmt_1137_PhiAck/phi_stmt_1145_ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(237)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(237)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(237) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1145_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1145_ack_3159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1145_ack_0, ack => convolution3D_CP_1120_elements(237)); -- 
    -- CP-element group 238:  join  fork  transition  place  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	236 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	136 
    -- CP-element group 238: 	139 
    -- CP-element group 238:  members (10) 
      -- CP-element group 238: 	 branch_block_stmt_435/merge_stmt_1137__exit__
      -- CP-element group 238: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181__entry__
      -- CP-element group 238: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/RPIPE_maxpool_input_pipe_1154_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/RPIPE_maxpool_input_pipe_1154_Sample/rr
      -- CP-element group 238: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/RPIPE_maxpool_input_pipe_1154_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/$entry
      -- CP-element group 238: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/type_cast_1158_Update/cr
      -- CP-element group 238: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/type_cast_1158_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_435/assign_stmt_1155_to_assign_stmt_1181/type_cast_1158_update_start_
      -- CP-element group 238: 	 branch_block_stmt_435/merge_stmt_1137_PhiAck/$exit
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(238)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(238)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(238) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:RPIPE_maxpool_input_pipe_1154_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1158_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    rr_2357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(238), ack => RPIPE_maxpool_input_pipe_1154_inst_req_0); -- 
    cr_2376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(238), ack => type_cast_1158_inst_req_1); -- 
    convolution3D_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(236) & convolution3D_CP_1120_elements(237);
      gj_convolution3D_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	140 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (2) 
      -- CP-element group 239: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/type_cast_1192/SplitProtocol/Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/type_cast_1192/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(239)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(239)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(239) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1192_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1192_inst_ack_0, ack => convolution3D_CP_1120_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	140 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (2) 
      -- CP-element group 240: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/type_cast_1192/SplitProtocol/Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/type_cast_1192/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(240)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(240)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(240) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1192_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1192_inst_ack_1, ack => convolution3D_CP_1120_elements(240)); -- 
    -- CP-element group 241:  join  transition  place  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (8) 
      -- CP-element group 241: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/$exit
      -- CP-element group 241: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/$exit
      -- CP-element group 241: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/$exit
      -- CP-element group 241: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/type_cast_1192/$exit
      -- CP-element group 241: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_sources/type_cast_1192/SplitProtocol/$exit
      -- CP-element group 241: 	 branch_block_stmt_435/forx_xbodyx_xi181_getRemainingElementsx_xexit188_PhiReq/phi_stmt_1189/phi_stmt_1189_req
      -- CP-element group 241: 	 branch_block_stmt_435/merge_stmt_1188_PhiReqMerge
      -- CP-element group 241: 	 branch_block_stmt_435/merge_stmt_1188_PhiAck/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(241)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(241)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(241) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1189_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1189_req_3189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1189_req_3189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(241), ack => phi_stmt_1189_req_0); -- 
    convolution3D_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(239) & convolution3D_CP_1120_elements(240);
      gj_convolution3D_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	142 
    -- CP-element group 242: 	143 
    -- CP-element group 242: 	145 
    -- CP-element group 242: 	147 
    -- CP-element group 242:  members (29) 
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_index_scale_1/$entry
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_index_resize_1/index_resize_req
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_index_resize_1/$exit
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_index_resize_1/$entry
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_index_computed_1
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_index_scaled_1
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_index_resize_1/index_resize_ack
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_index_resized_1
      -- CP-element group 242: 	 branch_block_stmt_435/merge_stmt_1188__exit__
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227__entry__
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_final_index_sum_regn_Update/req
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/addr_of_1222_update_start_
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/$entry
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_final_index_sum_regn_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Update/word_access_complete/word_0/cr
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Update/word_access_complete/word_0/$entry
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_final_index_sum_regn_Sample/req
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Update/word_access_complete/$entry
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_final_index_sum_regn_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_final_index_sum_regn_update_start
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_index_scale_1/scale_rename_ack
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_index_scale_1/scale_rename_req
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/ptr_deref_1225_update_start_
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/addr_of_1222_complete/req
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/array_obj_ref_1221_index_scale_1/$exit
      -- CP-element group 242: 	 branch_block_stmt_435/assign_stmt_1199_to_assign_stmt_1227/addr_of_1222_complete/$entry
      -- CP-element group 242: 	 branch_block_stmt_435/merge_stmt_1188_PhiAck/$exit
      -- CP-element group 242: 	 branch_block_stmt_435/merge_stmt_1188_PhiAck/phi_stmt_1189_ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(242)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(242)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(242) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1189_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_1221_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:ptr_deref_1225_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:array_obj_ref_1221_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:addr_of_1222_final_reg_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1189_ack_3194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1189_ack_0, ack => convolution3D_CP_1120_elements(242)); -- 
    req_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(242), ack => array_obj_ref_1221_index_offset_req_1); -- 
    cr_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(242), ack => ptr_deref_1225_store_0_req_1); -- 
    req_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(242), ack => array_obj_ref_1221_index_offset_req_0); -- 
    req_2444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(242), ack => addr_of_1222_final_reg_req_1); -- 
    -- CP-element group 243:  merge  fork  transition  place  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	130 
    -- CP-element group 243: 	148 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	149 
    -- CP-element group 243: 	150 
    -- CP-element group 243:  members (13) 
      -- CP-element group 243: 	 branch_block_stmt_435/call_stmt_1232/call_stmt_1232_Update/ccr
      -- CP-element group 243: 	 branch_block_stmt_435/merge_stmt_1229__exit__
      -- CP-element group 243: 	 branch_block_stmt_435/call_stmt_1232__entry__
      -- CP-element group 243: 	 branch_block_stmt_435/call_stmt_1232/call_stmt_1232_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_435/call_stmt_1232/call_stmt_1232_Sample/crr
      -- CP-element group 243: 	 branch_block_stmt_435/call_stmt_1232/call_stmt_1232_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_435/call_stmt_1232/call_stmt_1232_update_start_
      -- CP-element group 243: 	 branch_block_stmt_435/call_stmt_1232/call_stmt_1232_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_435/call_stmt_1232/$entry
      -- CP-element group 243: 	 branch_block_stmt_435/merge_stmt_1229_PhiReqMerge
      -- CP-element group 243: 	 branch_block_stmt_435/merge_stmt_1229_PhiAck/$entry
      -- CP-element group 243: 	 branch_block_stmt_435/merge_stmt_1229_PhiAck/$exit
      -- CP-element group 243: 	 branch_block_stmt_435/merge_stmt_1229_PhiAck/dummy
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(243)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(243)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(243) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1232_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1232_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ccr_2511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(243), ack => call_stmt_1232_call_req_1); -- 
    crr_2506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(243), ack => call_stmt_1232_call_req_0); -- 
    convolution3D_CP_1120_elements(243) <= OrReduce(convolution3D_CP_1120_elements(130) & convolution3D_CP_1120_elements(148));
    -- CP-element group 244:  transition  output  delay-element  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	161 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	248 
    -- CP-element group 244:  members (5) 
      -- CP-element group 244: 	 branch_block_stmt_435/ifx_xend107_whilex_xbody_PhiReq/$exit
      -- CP-element group 244: 	 branch_block_stmt_435/ifx_xend107_whilex_xbody_PhiReq/phi_stmt_1299/$exit
      -- CP-element group 244: 	 branch_block_stmt_435/ifx_xend107_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/$exit
      -- CP-element group 244: 	 branch_block_stmt_435/ifx_xend107_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/type_cast_1305_konst_delay_trans
      -- CP-element group 244: 	 branch_block_stmt_435/ifx_xend107_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(244)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(244)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(244) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1299_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1299_req_3216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1299_req_3216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(244), ack => phi_stmt_1299_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(244) is a control-delay.
    cp_element_244_delay: control_delay_element  generic map(name => " 244_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(161), ack => convolution3D_CP_1120_elements(244), clk => clk, reset =>reset);
    -- CP-element group 245:  transition  input  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	173 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (2) 
      -- CP-element group 245: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/type_cast_1302/SplitProtocol/Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/type_cast_1302/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(245)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(245)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(245) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1302_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1302_inst_ack_0, ack => convolution3D_CP_1120_elements(245)); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	173 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (2) 
      -- CP-element group 246: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/type_cast_1302/SplitProtocol/Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/type_cast_1302/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(246)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(246)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(246) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1302_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1302_inst_ack_1, ack => convolution3D_CP_1120_elements(246)); -- 
    -- CP-element group 247:  join  transition  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- CP-element group 247: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/$exit
      -- CP-element group 247: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/$exit
      -- CP-element group 247: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/type_cast_1302/$exit
      -- CP-element group 247: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_sources/type_cast_1302/SplitProtocol/$exit
      -- CP-element group 247: 	 branch_block_stmt_435/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1299/phi_stmt_1299_req
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(247)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(247)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(247) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1299_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1299_req_3242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1299_req_3242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(247), ack => phi_stmt_1299_req_0); -- 
    convolution3D_cp_element_group_247: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_247"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(245) & convolution3D_CP_1120_elements(246);
      gj_convolution3D_cp_element_group_247 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(247), clk => clk, reset => reset); --
    end block;
    -- CP-element group 248:  merge  transition  place  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	244 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (2) 
      -- CP-element group 248: 	 branch_block_stmt_435/merge_stmt_1298_PhiReqMerge
      -- CP-element group 248: 	 branch_block_stmt_435/merge_stmt_1298_PhiAck/$entry
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(248)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(248)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(248) fired."); 
        -- 
      end if; --
    end process; 
    convolution3D_CP_1120_elements(248) <= OrReduce(convolution3D_CP_1120_elements(244) & convolution3D_CP_1120_elements(247));
    -- CP-element group 249:  fork  transition  place  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	162 
    -- CP-element group 249: 	163 
    -- CP-element group 249: 	164 
    -- CP-element group 249: 	165 
    -- CP-element group 249: 	168 
    -- CP-element group 249: 	169 
    -- CP-element group 249: 	170 
    -- CP-element group 249:  members (26) 
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1319_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1319_update_start_
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1327_Update/ccr
      -- CP-element group 249: 	 branch_block_stmt_435/merge_stmt_1298__exit__
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345__entry__
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1334_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1327_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1319_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1327_update_start_
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/$entry
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1323_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1334_Update/ccr
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1323_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1334_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1323_Sample/rr
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1334_Sample/crr
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1323_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1323_update_start_
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1334_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1323_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1319_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1319_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/call_stmt_1334_update_start_
      -- CP-element group 249: 	 branch_block_stmt_435/assign_stmt_1311_to_assign_stmt_1345/type_cast_1319_Sample/rr
      -- CP-element group 249: 	 branch_block_stmt_435/merge_stmt_1298_PhiAck/$exit
      -- CP-element group 249: 	 branch_block_stmt_435/merge_stmt_1298_PhiAck/phi_stmt_1299_ack
      -- 
    -- logger for CP element group convolution3D_CP_1120_elements(249)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolution3D_CP_1120_elements(249)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:convolution3D_CP_1120_elements(249) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:phi_stmt_1299_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1327_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1323_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1334_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1323_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:call_stmt_1334_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1319_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolution3D:CP:type_cast_1319_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1299_ack_3247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1299_ack_0, ack => convolution3D_CP_1120_elements(249)); -- 
    ccr_2629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(249), ack => call_stmt_1327_call_req_1); -- 
    cr_2615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(249), ack => type_cast_1323_inst_req_1); -- 
    ccr_2643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(249), ack => call_stmt_1334_call_req_1); -- 
    rr_2610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(249), ack => type_cast_1323_inst_req_0); -- 
    crr_2638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(249), ack => call_stmt_1334_call_req_0); -- 
    cr_2601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(249), ack => type_cast_1319_inst_req_1); -- 
    rr_2596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(249), ack => type_cast_1319_inst_req_0); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1081_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_495_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_692_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_875_wire : std_logic_vector(63 downto 0);
    signal R_indvar240_975_resized : std_logic_vector(13 downto 0);
    signal R_indvar240_975_scaled : std_logic_vector(13 downto 0);
    signal R_indvar256_586_resized : std_logic_vector(13 downto 0);
    signal R_indvar256_586_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_826_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_826_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1220_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1220_scaled : std_logic_vector(13 downto 0);
    signal add30_632 : std_logic_vector(63 downto 0);
    signal add36_650 : std_logic_vector(63 downto 0);
    signal add75_1003 : std_logic_vector(63 downto 0);
    signal add81_1021 : std_logic_vector(63 downto 0);
    signal add87_1039 : std_logic_vector(63 downto 0);
    signal add_614 : std_logic_vector(63 downto 0);
    signal addx_xi177_1164 : std_logic_vector(63 downto 0);
    signal addx_xi_770 : std_logic_vector(63 downto 0);
    signal and97_1099 : std_logic_vector(63 downto 0);
    signal and_710 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1221_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1221_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1221_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1221_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1221_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1221_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_587_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_587_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_587_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_587_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_587_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_587_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_827_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_827_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_827_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_827_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_827_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_827_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_976_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_976_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_976_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_976_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_976_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_976_root_address : std_logic_vector(13 downto 0);
    signal arrayidx106_1223 : std_logic_vector(31 downto 0);
    signal arrayidx47_829 : std_logic_vector(31 downto 0);
    signal arrayidx91_978 : std_logic_vector(31 downto 0);
    signal arrayidx_589 : std_logic_vector(31 downto 0);
    signal call109_1232 : std_logic_vector(63 downto 0);
    signal call164_1360 : std_logic_vector(63 downto 0);
    signal call19_592 : std_logic_vector(15 downto 0);
    signal call1_441 : std_logic_vector(15 downto 0);
    signal call22_605 : std_logic_vector(15 downto 0);
    signal call27_623 : std_logic_vector(15 downto 0);
    signal call2_444 : std_logic_vector(15 downto 0);
    signal call33_641 : std_logic_vector(15 downto 0);
    signal call3_447 : std_logic_vector(15 downto 0);
    signal call4_450 : std_logic_vector(15 downto 0);
    signal call5_453 : std_logic_vector(15 downto 0);
    signal call68_981 : std_logic_vector(15 downto 0);
    signal call6_456 : std_logic_vector(15 downto 0);
    signal call72_994 : std_logic_vector(15 downto 0);
    signal call78_1012 : std_logic_vector(15 downto 0);
    signal call7_459 : std_logic_vector(15 downto 0);
    signal call84_1030 : std_logic_vector(15 downto 0);
    signal call_438 : std_logic_vector(15 downto 0);
    signal callx_xi175_1155 : std_logic_vector(15 downto 0);
    signal callx_xi_761 : std_logic_vector(15 downto 0);
    signal cmp195_503 : std_logic_vector(0 downto 0);
    signal cmp65191_883 : std_logic_vector(0 downto 0);
    signal conv110_1357 : std_logic_vector(63 downto 0);
    signal conv11_471 : std_logic_vector(63 downto 0);
    signal conv135_1320 : std_logic_vector(63 downto 0);
    signal conv13_497 : std_logic_vector(63 downto 0);
    signal conv141_1324 : std_logic_vector(63 downto 0);
    signal conv165_1365 : std_logic_vector(63 downto 0);
    signal conv20_596 : std_logic_vector(63 downto 0);
    signal conv24_609 : std_logic_vector(63 downto 0);
    signal conv29_627 : std_logic_vector(63 downto 0);
    signal conv35_645 : std_logic_vector(63 downto 0);
    signal conv51_839 : std_logic_vector(63 downto 0);
    signal conv54_843 : std_logic_vector(63 downto 0);
    signal conv57_847 : std_logic_vector(63 downto 0);
    signal conv59_877 : std_logic_vector(63 downto 0);
    signal conv5x_xi176_1159 : std_logic_vector(63 downto 0);
    signal conv5x_xi_765 : std_logic_vector(63 downto 0);
    signal conv69_985 : std_logic_vector(63 downto 0);
    signal conv74_998 : std_logic_vector(63 downto 0);
    signal conv80_1016 : std_logic_vector(63 downto 0);
    signal conv86_1034 : std_logic_vector(63 downto 0);
    signal conv9_467 : std_logic_vector(63 downto 0);
    signal conv_463 : std_logic_vector(63 downto 0);
    signal elementx_x015x_xi174_1145 : std_logic_vector(63 downto 0);
    signal elementx_x015x_xi_751 : std_logic_vector(63 downto 0);
    signal exitcond26_1054 : std_logic_vector(0 downto 0);
    signal exitcond2_787 : std_logic_vector(0 downto 0);
    signal exitcond37_665 : std_logic_vector(0 downto 0);
    signal exitcond7_1345 : std_logic_vector(0 downto 0);
    signal exitcond_1181 : std_logic_vector(0 downto 0);
    signal iNsTr_38_805 : std_logic_vector(63 downto 0);
    signal iNsTr_52_1199 : std_logic_vector(63 downto 0);
    signal incx_xi179_1176 : std_logic_vector(15 downto 0);
    signal incx_xi_782 : std_logic_vector(15 downto 0);
    signal indvar240_964 : std_logic_vector(63 downto 0);
    signal indvar256_575 : std_logic_vector(63 downto 0);
    signal indvar_1299 : std_logic_vector(31 downto 0);
    signal indvarx_xnext241_1049 : std_logic_vector(63 downto 0);
    signal indvarx_xnext257_660 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1340 : std_logic_vector(31 downto 0);
    signal ix_x0x_xlcssa_697 : std_logic_vector(63 downto 0);
    signal ix_x1x_xlcssa_1086 : std_logic_vector(63 downto 0);
    signal mul116_1238 : std_logic_vector(15 downto 0);
    signal mul129_1243 : std_logic_vector(15 downto 0);
    signal mul12_481 : std_logic_vector(63 downto 0);
    signal mul134_1311 : std_logic_vector(31 downto 0);
    signal mul140_1316 : std_logic_vector(31 downto 0);
    signal mul52_852 : std_logic_vector(63 downto 0);
    signal mul55_857 : std_logic_vector(63 downto 0);
    signal mul58_862 : std_logic_vector(63 downto 0);
    signal mul_476 : std_logic_vector(63 downto 0);
    signal mulx_xi185_1205 : std_logic_vector(63 downto 0);
    signal mulx_xi_811 : std_logic_vector(63 downto 0);
    signal nx_x016x_xi173_1138 : std_logic_vector(15 downto 0);
    signal nx_x016x_xi_744 : std_logic_vector(15 downto 0);
    signal phitmp199_1083 : std_logic_vector(63 downto 0);
    signal phitmp_694 : std_logic_vector(63 downto 0);
    signal ptr_deref_1041_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1041_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1041_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1041_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1041_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1041_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1225_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1225_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1225_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1225_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1225_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1225_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_652_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_652_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_652_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_652_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_652_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_652_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_831_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_831_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_831_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_831_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_831_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_831_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext171_868 : std_logic_vector(63 downto 0);
    signal sext_487 : std_logic_vector(63 downto 0);
    signal sh_promx_xi186_1211 : std_logic_vector(63 downto 0);
    signal sh_promx_xi_817 : std_logic_vector(63 downto 0);
    signal shl12x_xi187_1216 : std_logic_vector(63 downto 0);
    signal shl12x_xi_822 : std_logic_vector(63 downto 0);
    signal shl26_620 : std_logic_vector(63 downto 0);
    signal shl32_638 : std_logic_vector(63 downto 0);
    signal shl71_991 : std_logic_vector(63 downto 0);
    signal shl77_1009 : std_logic_vector(63 downto 0);
    signal shl83_1027 : std_logic_vector(63 downto 0);
    signal shl_602 : std_logic_vector(63 downto 0);
    signal shlx_xi178_1170 : std_logic_vector(63 downto 0);
    signal shlx_xi178x_xlcssa_1189 : std_logic_vector(63 downto 0);
    signal shlx_xi_776 : std_logic_vector(63 downto 0);
    signal shlx_xix_xlcssa_795 : std_logic_vector(63 downto 0);
    signal sub149_1262 : std_logic_vector(15 downto 0);
    signal sub169_1370 : std_logic_vector(63 downto 0);
    signal sub_1256 : std_logic_vector(15 downto 0);
    signal tmp10_1291 : std_logic_vector(31 downto 0);
    signal tmp11_1296 : std_logic_vector(31 downto 0);
    signal tmp14_906 : std_logic_vector(63 downto 0);
    signal tmp15_910 : std_logic_vector(63 downto 0);
    signal tmp16_915 : std_logic_vector(63 downto 0);
    signal tmp17_919 : std_logic_vector(63 downto 0);
    signal tmp18_924 : std_logic_vector(63 downto 0);
    signal tmp19_928 : std_logic_vector(63 downto 0);
    signal tmp1_741 : std_logic_vector(15 downto 0);
    signal tmp201_728 : std_logic_vector(15 downto 0);
    signal tmp203_733 : std_logic_vector(15 downto 0);
    signal tmp208_1117 : std_logic_vector(15 downto 0);
    signal tmp20_933 : std_logic_vector(63 downto 0);
    signal tmp210_1122 : std_logic_vector(15 downto 0);
    signal tmp212_1127 : std_logic_vector(15 downto 0);
    signal tmp216_1268 : std_logic_vector(15 downto 0);
    signal tmp21_937 : std_logic_vector(31 downto 0);
    signal tmp22_942 : std_logic_vector(63 downto 0);
    signal tmp235_896 : std_logic_vector(63 downto 0);
    signal tmp236_902 : std_logic_vector(0 downto 0);
    signal tmp237_1074 : std_logic_vector(63 downto 0);
    signal tmp23_948 : std_logic_vector(63 downto 0);
    signal tmp24_954 : std_logic_vector(0 downto 0);
    signal tmp250_516 : std_logic_vector(63 downto 0);
    signal tmp251_522 : std_logic_vector(0 downto 0);
    signal tmp253_685 : std_logic_vector(63 downto 0);
    signal tmp27_526 : std_logic_vector(63 downto 0);
    signal tmp28_530 : std_logic_vector(63 downto 0);
    signal tmp29_535 : std_logic_vector(63 downto 0);
    signal tmp30_539 : std_logic_vector(63 downto 0);
    signal tmp31_544 : std_logic_vector(63 downto 0);
    signal tmp32_548 : std_logic_vector(31 downto 0);
    signal tmp33_553 : std_logic_vector(63 downto 0);
    signal tmp34_559 : std_logic_vector(63 downto 0);
    signal tmp35_565 : std_logic_vector(0 downto 0);
    signal tmp3_1131 : std_logic_vector(1 downto 0);
    signal tmp4_1135 : std_logic_vector(15 downto 0);
    signal tmp5_1272 : std_logic_vector(31 downto 0);
    signal tmp6_1278 : std_logic_vector(31 downto 0);
    signal tmp8_1282 : std_logic_vector(31 downto 0);
    signal tmp9_1287 : std_logic_vector(15 downto 0);
    signal tmp_737 : std_logic_vector(1 downto 0);
    signal tobool98_1105 : std_logic_vector(0 downto 0);
    signal tobool_716 : std_logic_vector(0 downto 0);
    signal type_cast_1007_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1025_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1047_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1066_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1072_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1077_wire : std_logic_vector(63 downto 0);
    signal type_cast_1080_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1089_wire : std_logic_vector(63 downto 0);
    signal type_cast_1092_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1097_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1103_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1141_wire : std_logic_vector(15 downto 0);
    signal type_cast_1144_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1148_wire : std_logic_vector(63 downto 0);
    signal type_cast_1151_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1168_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1174_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1192_wire : std_logic_vector(63 downto 0);
    signal type_cast_1197_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1203_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1209_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1249_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1254_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1260_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1266_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1276_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1302_wire : std_logic_vector(31 downto 0);
    signal type_cast_1305_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1338_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1355_wire : std_logic_vector(63 downto 0);
    signal type_cast_1363_wire : std_logic_vector(63 downto 0);
    signal type_cast_485_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_491_wire : std_logic_vector(63 downto 0);
    signal type_cast_494_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_501_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_514_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_520_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_551_wire : std_logic_vector(63 downto 0);
    signal type_cast_557_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_563_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_570_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_579_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_581_wire : std_logic_vector(63 downto 0);
    signal type_cast_600_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_618_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_636_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_658_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_677_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_683_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_688_wire : std_logic_vector(63 downto 0);
    signal type_cast_691_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_700_wire : std_logic_vector(63 downto 0);
    signal type_cast_703_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_708_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_714_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_747_wire : std_logic_vector(15 downto 0);
    signal type_cast_750_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_754_wire : std_logic_vector(63 downto 0);
    signal type_cast_757_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_774_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_780_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_798_wire : std_logic_vector(63 downto 0);
    signal type_cast_803_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_809_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_815_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_866_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_871_wire : std_logic_vector(63 downto 0);
    signal type_cast_874_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_881_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_894_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_900_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_940_wire : std_logic_vector(63 downto 0);
    signal type_cast_946_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_952_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_959_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_968_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_970_wire : std_logic_vector(63 downto 0);
    signal type_cast_989_wire_constant : std_logic_vector(63 downto 0);
    signal umax252_679 : std_logic_vector(63 downto 0);
    signal umax25_961 : std_logic_vector(63 downto 0);
    signal umax36_572 : std_logic_vector(63 downto 0);
    signal umax_1068 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1221_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1221_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1221_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1221_resized_base_address <= "00000000000000";
    array_obj_ref_587_constant_part_of_offset <= "00000000000000";
    array_obj_ref_587_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_587_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_587_resized_base_address <= "00000000000000";
    array_obj_ref_827_constant_part_of_offset <= "00000000000000";
    array_obj_ref_827_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_827_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_827_resized_base_address <= "00000000000000";
    array_obj_ref_976_constant_part_of_offset <= "00000000000000";
    array_obj_ref_976_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_976_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_976_resized_base_address <= "00000000000000";
    ptr_deref_1041_word_offset_0 <= "00000000000000";
    ptr_deref_1225_word_offset_0 <= "00000000000000";
    ptr_deref_652_word_offset_0 <= "00000000000000";
    ptr_deref_831_word_offset_0 <= "00000000000000";
    type_cast_1007_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1025_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1047_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1066_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1072_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1080_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1092_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1097_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1103_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1144_wire_constant <= "0000000000000000";
    type_cast_1151_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1168_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1174_wire_constant <= "0000000000000001";
    type_cast_1197_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1203_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1209_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1249_wire_constant <= "0000000100101100";
    type_cast_1254_wire_constant <= "1111111111111111";
    type_cast_1260_wire_constant <= "1111111111111111";
    type_cast_1266_wire_constant <= "1111111111111111";
    type_cast_1276_wire_constant <= "00000000000000000000000000000001";
    type_cast_1305_wire_constant <= "00000000000000000000000000000000";
    type_cast_1338_wire_constant <= "00000000000000000000000000000001";
    type_cast_485_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_494_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_501_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_514_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_520_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_557_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_563_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_570_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_579_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_600_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_618_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_636_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_658_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_677_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_683_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_691_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_703_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_708_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_714_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_750_wire_constant <= "0000000000000000";
    type_cast_757_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_774_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_780_wire_constant <= "0000000000000001";
    type_cast_803_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_809_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_815_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_866_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_874_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_881_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_894_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_900_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_946_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_952_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_959_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_968_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_989_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    -- logger for phi phi_stmt_1086
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1086_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_1086:input-0 type_cast_1089_wire= " & Convert_SLV_To_Hex_String(type_cast_1089_wire));
          --
        end if;
        if phi_stmt_1086_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_1086:input-1 type_cast_1092_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1092_wire_constant));
          --
        end if;
        if phi_stmt_1086_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolution3D:DP:phi_stmt_1086:sample-completed");
          --
        end if;
        if phi_stmt_1086_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolution3D:DP:phi_stmt_1086:output ix_x1x_xlcssa_1086= " & Convert_SLV_To_Hex_String(ix_x1x_xlcssa_1086));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1086: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1089_wire & type_cast_1092_wire_constant;
      req <= phi_stmt_1086_req_0 & phi_stmt_1086_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1086",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1086_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_1086,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1086
    -- logger for phi phi_stmt_1138
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1138_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_1138:input-0 type_cast_1141_wire= " & Convert_SLV_To_Hex_String(type_cast_1141_wire));
          --
        end if;
        if phi_stmt_1138_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_1138:input-1 type_cast_1144_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1144_wire_constant));
          --
        end if;
        if phi_stmt_1138_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolution3D:DP:phi_stmt_1138:sample-completed");
          --
        end if;
        if phi_stmt_1138_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolution3D:DP:phi_stmt_1138:output nx_x016x_xi173_1138= " & Convert_SLV_To_Hex_String(nx_x016x_xi173_1138));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1138: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1141_wire & type_cast_1144_wire_constant;
      req <= phi_stmt_1138_req_0 & phi_stmt_1138_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1138",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1138_ack_0,
          idata => idata,
          odata => nx_x016x_xi173_1138,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1138
    -- logger for phi phi_stmt_1145
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1145_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_1145:input-0 type_cast_1148_wire= " & Convert_SLV_To_Hex_String(type_cast_1148_wire));
          --
        end if;
        if phi_stmt_1145_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_1145:input-1 type_cast_1151_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1151_wire_constant));
          --
        end if;
        if phi_stmt_1145_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolution3D:DP:phi_stmt_1145:sample-completed");
          --
        end if;
        if phi_stmt_1145_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolution3D:DP:phi_stmt_1145:output elementx_x015x_xi174_1145= " & Convert_SLV_To_Hex_String(elementx_x015x_xi174_1145));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1145: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1148_wire & type_cast_1151_wire_constant;
      req <= phi_stmt_1145_req_0 & phi_stmt_1145_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1145",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1145_ack_0,
          idata => idata,
          odata => elementx_x015x_xi174_1145,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1145
    -- logger for phi phi_stmt_1189
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1189_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_1189:input-0 type_cast_1192_wire= " & Convert_SLV_To_Hex_String(type_cast_1192_wire));
          --
        end if;
        if phi_stmt_1189_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolution3D:DP:phi_stmt_1189:sample-completed");
          --
        end if;
        if phi_stmt_1189_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolution3D:DP:phi_stmt_1189:output shlx_xi178x_xlcssa_1189= " & Convert_SLV_To_Hex_String(shlx_xi178x_xlcssa_1189));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1189: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1192_wire;
      req(0) <= phi_stmt_1189_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1189",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1189_ack_0,
          idata => idata,
          odata => shlx_xi178x_xlcssa_1189,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1189
    -- logger for phi phi_stmt_1299
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1299_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_1299:input-0 type_cast_1302_wire= " & Convert_SLV_To_Hex_String(type_cast_1302_wire));
          --
        end if;
        if phi_stmt_1299_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_1299:input-1 type_cast_1305_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1305_wire_constant));
          --
        end if;
        if phi_stmt_1299_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolution3D:DP:phi_stmt_1299:sample-completed");
          --
        end if;
        if phi_stmt_1299_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolution3D:DP:phi_stmt_1299:output indvar_1299= " & Convert_SLV_To_Hex_String(indvar_1299));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1299: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1302_wire & type_cast_1305_wire_constant;
      req <= phi_stmt_1299_req_0 & phi_stmt_1299_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1299",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1299_ack_0,
          idata => idata,
          odata => indvar_1299,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1299
    -- logger for phi phi_stmt_575
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_575_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_575:input-0 type_cast_579_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_579_wire_constant));
          --
        end if;
        if phi_stmt_575_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_575:input-1 type_cast_581_wire= " & Convert_SLV_To_Hex_String(type_cast_581_wire));
          --
        end if;
        if phi_stmt_575_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolution3D:DP:phi_stmt_575:sample-completed");
          --
        end if;
        if phi_stmt_575_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolution3D:DP:phi_stmt_575:output indvar256_575= " & Convert_SLV_To_Hex_String(indvar256_575));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_575: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_579_wire_constant & type_cast_581_wire;
      req <= phi_stmt_575_req_0 & phi_stmt_575_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_575",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_575_ack_0,
          idata => idata,
          odata => indvar256_575,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_575
    -- logger for phi phi_stmt_697
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_697_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_697:input-0 type_cast_700_wire= " & Convert_SLV_To_Hex_String(type_cast_700_wire));
          --
        end if;
        if phi_stmt_697_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_697:input-1 type_cast_703_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_703_wire_constant));
          --
        end if;
        if phi_stmt_697_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolution3D:DP:phi_stmt_697:sample-completed");
          --
        end if;
        if phi_stmt_697_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolution3D:DP:phi_stmt_697:output ix_x0x_xlcssa_697= " & Convert_SLV_To_Hex_String(ix_x0x_xlcssa_697));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_697: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_700_wire & type_cast_703_wire_constant;
      req <= phi_stmt_697_req_0 & phi_stmt_697_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_697",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_697_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_697,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_697
    -- logger for phi phi_stmt_744
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_744_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_744:input-0 type_cast_747_wire= " & Convert_SLV_To_Hex_String(type_cast_747_wire));
          --
        end if;
        if phi_stmt_744_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_744:input-1 type_cast_750_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_750_wire_constant));
          --
        end if;
        if phi_stmt_744_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolution3D:DP:phi_stmt_744:sample-completed");
          --
        end if;
        if phi_stmt_744_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolution3D:DP:phi_stmt_744:output nx_x016x_xi_744= " & Convert_SLV_To_Hex_String(nx_x016x_xi_744));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_744: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_747_wire & type_cast_750_wire_constant;
      req <= phi_stmt_744_req_0 & phi_stmt_744_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_744",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_744_ack_0,
          idata => idata,
          odata => nx_x016x_xi_744,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_744
    -- logger for phi phi_stmt_751
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_751_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_751:input-0 type_cast_754_wire= " & Convert_SLV_To_Hex_String(type_cast_754_wire));
          --
        end if;
        if phi_stmt_751_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_751:input-1 type_cast_757_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_757_wire_constant));
          --
        end if;
        if phi_stmt_751_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolution3D:DP:phi_stmt_751:sample-completed");
          --
        end if;
        if phi_stmt_751_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolution3D:DP:phi_stmt_751:output elementx_x015x_xi_751= " & Convert_SLV_To_Hex_String(elementx_x015x_xi_751));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_751: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_754_wire & type_cast_757_wire_constant;
      req <= phi_stmt_751_req_0 & phi_stmt_751_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_751",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_751_ack_0,
          idata => idata,
          odata => elementx_x015x_xi_751,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_751
    -- logger for phi phi_stmt_795
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_795_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_795:input-0 type_cast_798_wire= " & Convert_SLV_To_Hex_String(type_cast_798_wire));
          --
        end if;
        if phi_stmt_795_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolution3D:DP:phi_stmt_795:sample-completed");
          --
        end if;
        if phi_stmt_795_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolution3D:DP:phi_stmt_795:output shlx_xix_xlcssa_795= " & Convert_SLV_To_Hex_String(shlx_xix_xlcssa_795));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_795: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_798_wire;
      req(0) <= phi_stmt_795_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_795",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_795_ack_0,
          idata => idata,
          odata => shlx_xix_xlcssa_795,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_795
    -- logger for phi phi_stmt_964
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_964_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_964:input-0 type_cast_968_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_968_wire_constant));
          --
        end if;
        if phi_stmt_964_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolution3D:DP:phi_stmt_964:input-1 type_cast_970_wire= " & Convert_SLV_To_Hex_String(type_cast_970_wire));
          --
        end if;
        if phi_stmt_964_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolution3D:DP:phi_stmt_964:sample-completed");
          --
        end if;
        if phi_stmt_964_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolution3D:DP:phi_stmt_964:output indvar240_964= " & Convert_SLV_To_Hex_String(indvar240_964));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_964: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_968_wire_constant & type_cast_970_wire;
      req <= phi_stmt_964_req_0 & phi_stmt_964_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_964",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_964_ack_0,
          idata => idata,
          odata => indvar240_964,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_964
    -- logger for split-operator MUX_1067_inst flow-through 
    process(umax_1068) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUX_1067_inst:flowthrough inputs: " & " tmp236_902 = "& Convert_SLV_To_Hex_String(tmp236_902) & " tmp235_896 = "& Convert_SLV_To_Hex_String(tmp235_896) & " type_cast_1066_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1066_wire_constant) & " outputs:" & " umax_1068= "  & Convert_SLV_To_Hex_String(umax_1068));
      --
    end process; 
    -- flow-through select operator MUX_1067_inst
    umax_1068 <= tmp235_896 when (tmp236_902(0) /=  '0') else type_cast_1066_wire_constant;
    -- logger for split-operator MUX_571_inst flow-through 
    process(umax36_572) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUX_571_inst:flowthrough inputs: " & " tmp35_565 = "& Convert_SLV_To_Hex_String(tmp35_565) & " tmp34_559 = "& Convert_SLV_To_Hex_String(tmp34_559) & " type_cast_570_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_570_wire_constant) & " outputs:" & " umax36_572= "  & Convert_SLV_To_Hex_String(umax36_572));
      --
    end process; 
    -- flow-through select operator MUX_571_inst
    umax36_572 <= tmp34_559 when (tmp35_565(0) /=  '0') else type_cast_570_wire_constant;
    -- logger for split-operator MUX_678_inst flow-through 
    process(umax252_679) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUX_678_inst:flowthrough inputs: " & " tmp251_522 = "& Convert_SLV_To_Hex_String(tmp251_522) & " tmp250_516 = "& Convert_SLV_To_Hex_String(tmp250_516) & " type_cast_677_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_677_wire_constant) & " outputs:" & " umax252_679= "  & Convert_SLV_To_Hex_String(umax252_679));
      --
    end process; 
    -- flow-through select operator MUX_678_inst
    umax252_679 <= tmp250_516 when (tmp251_522(0) /=  '0') else type_cast_677_wire_constant;
    -- logger for split-operator MUX_960_inst flow-through 
    process(umax25_961) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUX_960_inst:flowthrough inputs: " & " tmp24_954 = "& Convert_SLV_To_Hex_String(tmp24_954) & " tmp23_948 = "& Convert_SLV_To_Hex_String(tmp23_948) & " type_cast_959_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_959_wire_constant) & " outputs:" & " umax25_961= "  & Convert_SLV_To_Hex_String(umax25_961));
      --
    end process; 
    -- flow-through select operator MUX_960_inst
    umax25_961 <= tmp23_948 when (tmp24_954(0) /=  '0') else type_cast_959_wire_constant;
    -- logger for split-operator addr_of_1222_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_1222_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:addr_of_1222_final_reg:started:   inputs: " & " array_obj_ref_1221_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1221_root_address));
          --
        end if; 
        if addr_of_1222_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:addr_of_1222_final_reg:finished:  outputs: " & " arrayidx106_1223= "  & Convert_SLV_To_Hex_String(arrayidx106_1223));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_1222_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1222_final_reg_req_0;
      addr_of_1222_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1222_final_reg_req_1;
      addr_of_1222_final_reg_ack_1<= rack(0);
      addr_of_1222_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1222_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1221_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx106_1223,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_588_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_588_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:addr_of_588_final_reg:started:   inputs: " & " array_obj_ref_587_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_587_root_address));
          --
        end if; 
        if addr_of_588_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:addr_of_588_final_reg:finished:  outputs: " & " arrayidx_589= "  & Convert_SLV_To_Hex_String(arrayidx_589));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_588_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_588_final_reg_req_0;
      addr_of_588_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_588_final_reg_req_1;
      addr_of_588_final_reg_ack_1<= rack(0);
      addr_of_588_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_588_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_587_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_589,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_828_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_828_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:addr_of_828_final_reg:started:   inputs: " & " array_obj_ref_827_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_827_root_address));
          --
        end if; 
        if addr_of_828_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:addr_of_828_final_reg:finished:  outputs: " & " arrayidx47_829= "  & Convert_SLV_To_Hex_String(arrayidx47_829));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_828_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_828_final_reg_req_0;
      addr_of_828_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_828_final_reg_req_1;
      addr_of_828_final_reg_ack_1<= rack(0);
      addr_of_828_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_828_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_827_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx47_829,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_977_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_977_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:addr_of_977_final_reg:started:   inputs: " & " array_obj_ref_976_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_976_root_address));
          --
        end if; 
        if addr_of_977_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:addr_of_977_final_reg:finished:  outputs: " & " arrayidx91_978= "  & Convert_SLV_To_Hex_String(arrayidx91_978));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_977_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_977_final_reg_req_0;
      addr_of_977_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_977_final_reg_req_1;
      addr_of_977_final_reg_ack_1<= rack(0);
      addr_of_977_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_977_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_976_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx91_978,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1015_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1015_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1015_inst:started:   inputs: " & " call78_1012 = "& Convert_SLV_To_Hex_String(call78_1012));
          --
        end if; 
        if type_cast_1015_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1015_inst:finished:  outputs: " & " conv80_1016= "  & Convert_SLV_To_Hex_String(conv80_1016));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1015_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1015_inst_req_0;
      type_cast_1015_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1015_inst_req_1;
      type_cast_1015_inst_ack_1<= rack(0);
      type_cast_1015_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1015_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call78_1012,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_1016,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1033_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1033_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1033_inst:started:   inputs: " & " call84_1030 = "& Convert_SLV_To_Hex_String(call84_1030));
          --
        end if; 
        if type_cast_1033_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1033_inst:finished:  outputs: " & " conv86_1034= "  & Convert_SLV_To_Hex_String(conv86_1034));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1033_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1033_inst_req_0;
      type_cast_1033_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1033_inst_req_1;
      type_cast_1033_inst_ack_1<= rack(0);
      type_cast_1033_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1033_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call84_1030,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_1034,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1077_inst flow-through 
    process(type_cast_1077_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1077_inst:flowthrough inputs: " & " tmp237_1074 = "& Convert_SLV_To_Hex_String(tmp237_1074) & " outputs:" & " type_cast_1077_wire= "  & Convert_SLV_To_Hex_String(type_cast_1077_wire));
      --
    end process; 
    -- interlock type_cast_1077_inst
    process(tmp237_1074) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp237_1074(63 downto 0);
      type_cast_1077_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1082_inst flow-through 
    process(phitmp199_1083) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1082_inst:flowthrough inputs: " & " ASHR_i64_i64_1081_wire = "& Convert_SLV_To_Hex_String(ASHR_i64_i64_1081_wire) & " outputs:" & " phitmp199_1083= "  & Convert_SLV_To_Hex_String(phitmp199_1083));
      --
    end process; 
    -- interlock type_cast_1082_inst
    process(ASHR_i64_i64_1081_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1081_wire(63 downto 0);
      phitmp199_1083 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1089_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1089_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1089_inst:started:   inputs: " & " phitmp199_1083 = "& Convert_SLV_To_Hex_String(phitmp199_1083));
          --
        end if; 
        if type_cast_1089_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1089_inst:finished:  outputs: " & " type_cast_1089_wire= "  & Convert_SLV_To_Hex_String(type_cast_1089_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1089_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1089_inst_req_0;
      type_cast_1089_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1089_inst_req_1;
      type_cast_1089_inst_ack_1<= rack(0);
      type_cast_1089_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1089_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp199_1083,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1089_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1130_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1130_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1130_inst:started:   inputs: " & " tmp212_1127 = "& Convert_SLV_To_Hex_String(tmp212_1127));
          --
        end if; 
        if type_cast_1130_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1130_inst:finished:  outputs: " & " tmp3_1131= "  & Convert_SLV_To_Hex_String(tmp3_1131));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1130_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1130_inst_req_0;
      type_cast_1130_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1130_inst_req_1;
      type_cast_1130_inst_ack_1<= rack(0);
      type_cast_1130_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1130_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp212_1127,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_1131,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1134_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1134_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1134_inst:started:   inputs: " & " tmp3_1131 = "& Convert_SLV_To_Hex_String(tmp3_1131));
          --
        end if; 
        if type_cast_1134_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1134_inst:finished:  outputs: " & " tmp4_1135= "  & Convert_SLV_To_Hex_String(tmp4_1135));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1134_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1134_inst_req_0;
      type_cast_1134_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1134_inst_req_1;
      type_cast_1134_inst_ack_1<= rack(0);
      type_cast_1134_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1134_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_1131,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp4_1135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1141_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1141_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1141_inst:started:   inputs: " & " incx_xi179_1176 = "& Convert_SLV_To_Hex_String(incx_xi179_1176));
          --
        end if; 
        if type_cast_1141_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1141_inst:finished:  outputs: " & " type_cast_1141_wire= "  & Convert_SLV_To_Hex_String(type_cast_1141_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1141_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1141_inst_req_0;
      type_cast_1141_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1141_inst_req_1;
      type_cast_1141_inst_ack_1<= rack(0);
      type_cast_1141_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1141_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => incx_xi179_1176,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1141_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1148_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1148_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1148_inst:started:   inputs: " & " shlx_xi178_1170 = "& Convert_SLV_To_Hex_String(shlx_xi178_1170));
          --
        end if; 
        if type_cast_1148_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1148_inst:finished:  outputs: " & " type_cast_1148_wire= "  & Convert_SLV_To_Hex_String(type_cast_1148_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1148_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1148_inst_req_0;
      type_cast_1148_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1148_inst_req_1;
      type_cast_1148_inst_ack_1<= rack(0);
      type_cast_1148_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1148_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shlx_xi178_1170,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1148_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1158_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1158_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1158_inst:started:   inputs: " & " callx_xi175_1155 = "& Convert_SLV_To_Hex_String(callx_xi175_1155));
          --
        end if; 
        if type_cast_1158_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1158_inst:finished:  outputs: " & " conv5x_xi176_1159= "  & Convert_SLV_To_Hex_String(conv5x_xi176_1159));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1158_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1158_inst_req_0;
      type_cast_1158_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1158_inst_req_1;
      type_cast_1158_inst_ack_1<= rack(0);
      type_cast_1158_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1158_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi175_1155,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi176_1159,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1192_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1192_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1192_inst:started:   inputs: " & " shlx_xi178_1170 = "& Convert_SLV_To_Hex_String(shlx_xi178_1170));
          --
        end if; 
        if type_cast_1192_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1192_inst:finished:  outputs: " & " type_cast_1192_wire= "  & Convert_SLV_To_Hex_String(type_cast_1192_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1192_inst_req_0;
      type_cast_1192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1192_inst_req_1;
      type_cast_1192_inst_ack_1<= rack(0);
      type_cast_1192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shlx_xi178_1170,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1192_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1271_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1271_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1271_inst:started:   inputs: " & " tmp216_1268 = "& Convert_SLV_To_Hex_String(tmp216_1268));
          --
        end if; 
        if type_cast_1271_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1271_inst:finished:  outputs: " & " tmp5_1272= "  & Convert_SLV_To_Hex_String(tmp5_1272));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1271_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1271_inst_req_0;
      type_cast_1271_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1271_inst_req_1;
      type_cast_1271_inst_ack_1<= rack(0);
      type_cast_1271_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1271_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp216_1268,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp5_1272,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1281_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1281_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1281_inst:started:   inputs: " & " call6_456 = "& Convert_SLV_To_Hex_String(call6_456));
          --
        end if; 
        if type_cast_1281_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1281_inst:finished:  outputs: " & " tmp8_1282= "  & Convert_SLV_To_Hex_String(tmp8_1282));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1281_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1281_inst_req_0;
      type_cast_1281_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1281_inst_req_1;
      type_cast_1281_inst_ack_1<= rack(0);
      type_cast_1281_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1281_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_456,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp8_1282,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1290_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1290_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1290_inst:started:   inputs: " & " tmp9_1287 = "& Convert_SLV_To_Hex_String(tmp9_1287));
          --
        end if; 
        if type_cast_1290_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1290_inst:finished:  outputs: " & " tmp10_1291= "  & Convert_SLV_To_Hex_String(tmp10_1291));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1290_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1290_inst_req_0;
      type_cast_1290_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1290_inst_req_1;
      type_cast_1290_inst_ack_1<= rack(0);
      type_cast_1290_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1290_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp9_1287,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp10_1291,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1302_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1302_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1302_inst:started:   inputs: " & " indvarx_xnext_1340 = "& Convert_SLV_To_Hex_String(indvarx_xnext_1340));
          --
        end if; 
        if type_cast_1302_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1302_inst:finished:  outputs: " & " type_cast_1302_wire= "  & Convert_SLV_To_Hex_String(type_cast_1302_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1302_inst_req_0;
      type_cast_1302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1302_inst_req_1;
      type_cast_1302_inst_ack_1<= rack(0);
      type_cast_1302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1340,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1302_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1319_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1319_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1319_inst:started:   inputs: " & " mul134_1311 = "& Convert_SLV_To_Hex_String(mul134_1311));
          --
        end if; 
        if type_cast_1319_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1319_inst:finished:  outputs: " & " conv135_1320= "  & Convert_SLV_To_Hex_String(conv135_1320));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1319_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1319_inst_req_0;
      type_cast_1319_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1319_inst_req_1;
      type_cast_1319_inst_ack_1<= rack(0);
      type_cast_1319_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1319_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul134_1311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv135_1320,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1323_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1323_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1323_inst:started:   inputs: " & " mul140_1316 = "& Convert_SLV_To_Hex_String(mul140_1316));
          --
        end if; 
        if type_cast_1323_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1323_inst:finished:  outputs: " & " conv141_1324= "  & Convert_SLV_To_Hex_String(conv141_1324));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1323_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1323_inst_req_0;
      type_cast_1323_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1323_inst_req_1;
      type_cast_1323_inst_ack_1<= rack(0);
      type_cast_1323_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1323_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul140_1316,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv141_1324,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1356_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1356_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1356_inst:started:   inputs: " & " type_cast_1355_wire = "& Convert_SLV_To_Hex_String(type_cast_1355_wire));
          --
        end if; 
        if type_cast_1356_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1356_inst:finished:  outputs: " & " conv110_1357= "  & Convert_SLV_To_Hex_String(conv110_1357));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1356_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1356_inst_req_0;
      type_cast_1356_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1356_inst_req_1;
      type_cast_1356_inst_ack_1<= rack(0);
      type_cast_1356_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1356_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1355_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_1357,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1364_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1364_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1364_inst:started:   inputs: " & " type_cast_1363_wire = "& Convert_SLV_To_Hex_String(type_cast_1363_wire));
          --
        end if; 
        if type_cast_1364_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1364_inst:finished:  outputs: " & " conv165_1365= "  & Convert_SLV_To_Hex_String(conv165_1365));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1364_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1364_inst_req_0;
      type_cast_1364_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1364_inst_req_1;
      type_cast_1364_inst_ack_1<= rack(0);
      type_cast_1364_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1364_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1363_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_1365,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_462_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_462_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_462_inst:started:   inputs: " & " call_438 = "& Convert_SLV_To_Hex_String(call_438));
          --
        end if; 
        if type_cast_462_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_462_inst:finished:  outputs: " & " conv_463= "  & Convert_SLV_To_Hex_String(conv_463));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_462_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_462_inst_req_0;
      type_cast_462_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_462_inst_req_1;
      type_cast_462_inst_ack_1<= rack(0);
      type_cast_462_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_462_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_438,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_463,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_466_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_466_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_466_inst:started:   inputs: " & " call1_441 = "& Convert_SLV_To_Hex_String(call1_441));
          --
        end if; 
        if type_cast_466_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_466_inst:finished:  outputs: " & " conv9_467= "  & Convert_SLV_To_Hex_String(conv9_467));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_466_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_466_inst_req_0;
      type_cast_466_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_466_inst_req_1;
      type_cast_466_inst_ack_1<= rack(0);
      type_cast_466_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_466_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_441,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_467,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_470_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_470_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_470_inst:started:   inputs: " & " call2_444 = "& Convert_SLV_To_Hex_String(call2_444));
          --
        end if; 
        if type_cast_470_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_470_inst:finished:  outputs: " & " conv11_471= "  & Convert_SLV_To_Hex_String(conv11_471));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_470_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_470_inst_req_0;
      type_cast_470_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_470_inst_req_1;
      type_cast_470_inst_ack_1<= rack(0);
      type_cast_470_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_470_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_444,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_471,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_491_inst flow-through 
    process(type_cast_491_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_491_inst:flowthrough inputs: " & " sext_487 = "& Convert_SLV_To_Hex_String(sext_487) & " outputs:" & " type_cast_491_wire= "  & Convert_SLV_To_Hex_String(type_cast_491_wire));
      --
    end process; 
    -- interlock type_cast_491_inst
    process(sext_487) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_487(63 downto 0);
      type_cast_491_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_496_inst flow-through 
    process(conv13_497) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_496_inst:flowthrough inputs: " & " ASHR_i64_i64_495_wire = "& Convert_SLV_To_Hex_String(ASHR_i64_i64_495_wire) & " outputs:" & " conv13_497= "  & Convert_SLV_To_Hex_String(conv13_497));
      --
    end process; 
    -- interlock type_cast_496_inst
    process(ASHR_i64_i64_495_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_495_wire(63 downto 0);
      conv13_497 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_525_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_525_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_525_inst:started:   inputs: " & " call1_441 = "& Convert_SLV_To_Hex_String(call1_441));
          --
        end if; 
        if type_cast_525_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_525_inst:finished:  outputs: " & " tmp27_526= "  & Convert_SLV_To_Hex_String(tmp27_526));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_525_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_525_inst_req_0;
      type_cast_525_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_525_inst_req_1;
      type_cast_525_inst_ack_1<= rack(0);
      type_cast_525_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_525_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_441,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp27_526,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_529_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_529_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_529_inst:started:   inputs: " & " call_438 = "& Convert_SLV_To_Hex_String(call_438));
          --
        end if; 
        if type_cast_529_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_529_inst:finished:  outputs: " & " tmp28_530= "  & Convert_SLV_To_Hex_String(tmp28_530));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_529_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_529_inst_req_0;
      type_cast_529_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_529_inst_req_1;
      type_cast_529_inst_ack_1<= rack(0);
      type_cast_529_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_529_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_438,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp28_530,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_538_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_538_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_538_inst:started:   inputs: " & " call2_444 = "& Convert_SLV_To_Hex_String(call2_444));
          --
        end if; 
        if type_cast_538_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_538_inst:finished:  outputs: " & " tmp30_539= "  & Convert_SLV_To_Hex_String(tmp30_539));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_538_inst_req_0;
      type_cast_538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_538_inst_req_1;
      type_cast_538_inst_ack_1<= rack(0);
      type_cast_538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_444,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp30_539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_547_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_547_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_547_inst:started:   inputs: " & " tmp31_544 = "& Convert_SLV_To_Hex_String(tmp31_544));
          --
        end if; 
        if type_cast_547_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_547_inst:finished:  outputs: " & " tmp32_548= "  & Convert_SLV_To_Hex_String(tmp32_548));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_547_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_547_inst_req_0;
      type_cast_547_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_547_inst_req_1;
      type_cast_547_inst_ack_1<= rack(0);
      type_cast_547_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_547_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp31_544,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp32_548,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_552_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_552_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_552_inst:started:   inputs: " & " type_cast_551_wire = "& Convert_SLV_To_Hex_String(type_cast_551_wire));
          --
        end if; 
        if type_cast_552_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_552_inst:finished:  outputs: " & " tmp33_553= "  & Convert_SLV_To_Hex_String(tmp33_553));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_552_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_552_inst_req_0;
      type_cast_552_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_552_inst_req_1;
      type_cast_552_inst_ack_1<= rack(0);
      type_cast_552_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_552_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_551_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp33_553,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_581_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_581_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_581_inst:started:   inputs: " & " indvarx_xnext257_660 = "& Convert_SLV_To_Hex_String(indvarx_xnext257_660));
          --
        end if; 
        if type_cast_581_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_581_inst:finished:  outputs: " & " type_cast_581_wire= "  & Convert_SLV_To_Hex_String(type_cast_581_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_581_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_581_inst_req_0;
      type_cast_581_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_581_inst_req_1;
      type_cast_581_inst_ack_1<= rack(0);
      type_cast_581_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_581_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext257_660,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_581_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_595_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_595_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_595_inst:started:   inputs: " & " call19_592 = "& Convert_SLV_To_Hex_String(call19_592));
          --
        end if; 
        if type_cast_595_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_595_inst:finished:  outputs: " & " conv20_596= "  & Convert_SLV_To_Hex_String(conv20_596));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_595_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_595_inst_req_0;
      type_cast_595_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_595_inst_req_1;
      type_cast_595_inst_ack_1<= rack(0);
      type_cast_595_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_595_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_592,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_596,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_608_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_608_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_608_inst:started:   inputs: " & " call22_605 = "& Convert_SLV_To_Hex_String(call22_605));
          --
        end if; 
        if type_cast_608_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_608_inst:finished:  outputs: " & " conv24_609= "  & Convert_SLV_To_Hex_String(conv24_609));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_608_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_608_inst_req_0;
      type_cast_608_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_608_inst_req_1;
      type_cast_608_inst_ack_1<= rack(0);
      type_cast_608_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_608_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_609,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_626_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_626_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_626_inst:started:   inputs: " & " call27_623 = "& Convert_SLV_To_Hex_String(call27_623));
          --
        end if; 
        if type_cast_626_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_626_inst:finished:  outputs: " & " conv29_627= "  & Convert_SLV_To_Hex_String(conv29_627));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_626_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_626_inst_req_0;
      type_cast_626_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_626_inst_req_1;
      type_cast_626_inst_ack_1<= rack(0);
      type_cast_626_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_626_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call27_623,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_627,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_644_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_644_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_644_inst:started:   inputs: " & " call33_641 = "& Convert_SLV_To_Hex_String(call33_641));
          --
        end if; 
        if type_cast_644_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_644_inst:finished:  outputs: " & " conv35_645= "  & Convert_SLV_To_Hex_String(conv35_645));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_644_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_644_inst_req_0;
      type_cast_644_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_644_inst_req_1;
      type_cast_644_inst_ack_1<= rack(0);
      type_cast_644_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_644_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call33_641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_645,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_688_inst flow-through 
    process(type_cast_688_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_688_inst:flowthrough inputs: " & " tmp253_685 = "& Convert_SLV_To_Hex_String(tmp253_685) & " outputs:" & " type_cast_688_wire= "  & Convert_SLV_To_Hex_String(type_cast_688_wire));
      --
    end process; 
    -- interlock type_cast_688_inst
    process(tmp253_685) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp253_685(63 downto 0);
      type_cast_688_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_693_inst flow-through 
    process(phitmp_694) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_693_inst:flowthrough inputs: " & " ASHR_i64_i64_692_wire = "& Convert_SLV_To_Hex_String(ASHR_i64_i64_692_wire) & " outputs:" & " phitmp_694= "  & Convert_SLV_To_Hex_String(phitmp_694));
      --
    end process; 
    -- interlock type_cast_693_inst
    process(ASHR_i64_i64_692_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_692_wire(63 downto 0);
      phitmp_694 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_700_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_700_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_700_inst:started:   inputs: " & " phitmp_694 = "& Convert_SLV_To_Hex_String(phitmp_694));
          --
        end if; 
        if type_cast_700_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_700_inst:finished:  outputs: " & " type_cast_700_wire= "  & Convert_SLV_To_Hex_String(type_cast_700_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_700_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_700_inst_req_0;
      type_cast_700_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_700_inst_req_1;
      type_cast_700_inst_ack_1<= rack(0);
      type_cast_700_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_700_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_694,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_700_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_736_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_736_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_736_inst:started:   inputs: " & " tmp203_733 = "& Convert_SLV_To_Hex_String(tmp203_733));
          --
        end if; 
        if type_cast_736_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_736_inst:finished:  outputs: " & " tmp_737= "  & Convert_SLV_To_Hex_String(tmp_737));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_736_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_736_inst_req_0;
      type_cast_736_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_736_inst_req_1;
      type_cast_736_inst_ack_1<= rack(0);
      type_cast_736_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_736_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp203_733,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp_737,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_740_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_740_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_740_inst:started:   inputs: " & " tmp_737 = "& Convert_SLV_To_Hex_String(tmp_737));
          --
        end if; 
        if type_cast_740_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_740_inst:finished:  outputs: " & " tmp1_741= "  & Convert_SLV_To_Hex_String(tmp1_741));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_740_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_740_inst_req_0;
      type_cast_740_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_740_inst_req_1;
      type_cast_740_inst_ack_1<= rack(0);
      type_cast_740_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_740_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_737,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_741,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_747_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_747_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_747_inst:started:   inputs: " & " incx_xi_782 = "& Convert_SLV_To_Hex_String(incx_xi_782));
          --
        end if; 
        if type_cast_747_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_747_inst:finished:  outputs: " & " type_cast_747_wire= "  & Convert_SLV_To_Hex_String(type_cast_747_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_747_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_747_inst_req_0;
      type_cast_747_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_747_inst_req_1;
      type_cast_747_inst_ack_1<= rack(0);
      type_cast_747_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_747_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => incx_xi_782,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_747_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_754_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_754_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_754_inst:started:   inputs: " & " shlx_xi_776 = "& Convert_SLV_To_Hex_String(shlx_xi_776));
          --
        end if; 
        if type_cast_754_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_754_inst:finished:  outputs: " & " type_cast_754_wire= "  & Convert_SLV_To_Hex_String(type_cast_754_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_754_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_754_inst_req_0;
      type_cast_754_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_754_inst_req_1;
      type_cast_754_inst_ack_1<= rack(0);
      type_cast_754_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_754_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shlx_xi_776,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_754_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_764_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_764_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_764_inst:started:   inputs: " & " callx_xi_761 = "& Convert_SLV_To_Hex_String(callx_xi_761));
          --
        end if; 
        if type_cast_764_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_764_inst:finished:  outputs: " & " conv5x_xi_765= "  & Convert_SLV_To_Hex_String(conv5x_xi_765));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_764_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_764_inst_req_0;
      type_cast_764_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_764_inst_req_1;
      type_cast_764_inst_ack_1<= rack(0);
      type_cast_764_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_764_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi_765,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_798_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_798_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_798_inst:started:   inputs: " & " shlx_xi_776 = "& Convert_SLV_To_Hex_String(shlx_xi_776));
          --
        end if; 
        if type_cast_798_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_798_inst:finished:  outputs: " & " type_cast_798_wire= "  & Convert_SLV_To_Hex_String(type_cast_798_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_798_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_798_inst_req_0;
      type_cast_798_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_798_inst_req_1;
      type_cast_798_inst_ack_1<= rack(0);
      type_cast_798_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_798_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shlx_xi_776,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_798_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_838_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_838_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_838_inst:started:   inputs: " & " call7_459 = "& Convert_SLV_To_Hex_String(call7_459));
          --
        end if; 
        if type_cast_838_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_838_inst:finished:  outputs: " & " conv51_839= "  & Convert_SLV_To_Hex_String(conv51_839));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_838_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_838_inst_req_0;
      type_cast_838_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_838_inst_req_1;
      type_cast_838_inst_ack_1<= rack(0);
      type_cast_838_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_838_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call7_459,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_839,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_842_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_842_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_842_inst:started:   inputs: " & " call6_456 = "& Convert_SLV_To_Hex_String(call6_456));
          --
        end if; 
        if type_cast_842_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_842_inst:finished:  outputs: " & " conv54_843= "  & Convert_SLV_To_Hex_String(conv54_843));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_842_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_842_inst_req_0;
      type_cast_842_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_842_inst_req_1;
      type_cast_842_inst_ack_1<= rack(0);
      type_cast_842_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_842_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_456,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv54_843,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_846_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_846_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_846_inst:started:   inputs: " & " call5_453 = "& Convert_SLV_To_Hex_String(call5_453));
          --
        end if; 
        if type_cast_846_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_846_inst:finished:  outputs: " & " conv57_847= "  & Convert_SLV_To_Hex_String(conv57_847));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_846_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_846_inst_req_0;
      type_cast_846_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_846_inst_req_1;
      type_cast_846_inst_ack_1<= rack(0);
      type_cast_846_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_846_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_453,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv57_847,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_871_inst flow-through 
    process(type_cast_871_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_871_inst:flowthrough inputs: " & " sext171_868 = "& Convert_SLV_To_Hex_String(sext171_868) & " outputs:" & " type_cast_871_wire= "  & Convert_SLV_To_Hex_String(type_cast_871_wire));
      --
    end process; 
    -- interlock type_cast_871_inst
    process(sext171_868) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext171_868(63 downto 0);
      type_cast_871_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_876_inst flow-through 
    process(conv59_877) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_876_inst:flowthrough inputs: " & " ASHR_i64_i64_875_wire = "& Convert_SLV_To_Hex_String(ASHR_i64_i64_875_wire) & " outputs:" & " conv59_877= "  & Convert_SLV_To_Hex_String(conv59_877));
      --
    end process; 
    -- interlock type_cast_876_inst
    process(ASHR_i64_i64_875_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_875_wire(63 downto 0);
      conv59_877 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_905_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_905_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_905_inst:started:   inputs: " & " call5_453 = "& Convert_SLV_To_Hex_String(call5_453));
          --
        end if; 
        if type_cast_905_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_905_inst:finished:  outputs: " & " tmp14_906= "  & Convert_SLV_To_Hex_String(tmp14_906));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_905_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_905_inst_req_0;
      type_cast_905_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_905_inst_req_1;
      type_cast_905_inst_ack_1<= rack(0);
      type_cast_905_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_905_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_453,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp14_906,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_909_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_909_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_909_inst:started:   inputs: " & " call2_444 = "& Convert_SLV_To_Hex_String(call2_444));
          --
        end if; 
        if type_cast_909_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_909_inst:finished:  outputs: " & " tmp15_910= "  & Convert_SLV_To_Hex_String(tmp15_910));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_909_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_909_inst_req_0;
      type_cast_909_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_909_inst_req_1;
      type_cast_909_inst_ack_1<= rack(0);
      type_cast_909_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_909_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_444,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_910,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_918_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_918_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_918_inst:started:   inputs: " & " call6_456 = "& Convert_SLV_To_Hex_String(call6_456));
          --
        end if; 
        if type_cast_918_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_918_inst:finished:  outputs: " & " tmp17_919= "  & Convert_SLV_To_Hex_String(tmp17_919));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_918_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_918_inst_req_0;
      type_cast_918_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_918_inst_req_1;
      type_cast_918_inst_ack_1<= rack(0);
      type_cast_918_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_918_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_456,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp17_919,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_927_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_927_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_927_inst:started:   inputs: " & " call7_459 = "& Convert_SLV_To_Hex_String(call7_459));
          --
        end if; 
        if type_cast_927_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_927_inst:finished:  outputs: " & " tmp19_928= "  & Convert_SLV_To_Hex_String(tmp19_928));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_927_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_927_inst_req_0;
      type_cast_927_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_927_inst_req_1;
      type_cast_927_inst_ack_1<= rack(0);
      type_cast_927_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_927_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call7_459,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp19_928,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_936_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_936_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_936_inst:started:   inputs: " & " tmp20_933 = "& Convert_SLV_To_Hex_String(tmp20_933));
          --
        end if; 
        if type_cast_936_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_936_inst:finished:  outputs: " & " tmp21_937= "  & Convert_SLV_To_Hex_String(tmp21_937));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_936_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_936_inst_req_0;
      type_cast_936_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_936_inst_req_1;
      type_cast_936_inst_ack_1<= rack(0);
      type_cast_936_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_936_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp20_933,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp21_937,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_941_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_941_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_941_inst:started:   inputs: " & " type_cast_940_wire = "& Convert_SLV_To_Hex_String(type_cast_940_wire));
          --
        end if; 
        if type_cast_941_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_941_inst:finished:  outputs: " & " tmp22_942= "  & Convert_SLV_To_Hex_String(tmp22_942));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_941_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_941_inst_req_0;
      type_cast_941_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_941_inst_req_1;
      type_cast_941_inst_ack_1<= rack(0);
      type_cast_941_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_941_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_940_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp22_942,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_970_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_970_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_970_inst:started:   inputs: " & " indvarx_xnext241_1049 = "& Convert_SLV_To_Hex_String(indvarx_xnext241_1049));
          --
        end if; 
        if type_cast_970_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_970_inst:finished:  outputs: " & " type_cast_970_wire= "  & Convert_SLV_To_Hex_String(type_cast_970_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_970_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_970_inst_req_0;
      type_cast_970_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_970_inst_req_1;
      type_cast_970_inst_ack_1<= rack(0);
      type_cast_970_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_970_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext241_1049,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_970_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_984_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_984_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_984_inst:started:   inputs: " & " call68_981 = "& Convert_SLV_To_Hex_String(call68_981));
          --
        end if; 
        if type_cast_984_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_984_inst:finished:  outputs: " & " conv69_985= "  & Convert_SLV_To_Hex_String(conv69_985));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_984_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_984_inst_req_0;
      type_cast_984_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_984_inst_req_1;
      type_cast_984_inst_ack_1<= rack(0);
      type_cast_984_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_984_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call68_981,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_985,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_997_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_997_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_997_inst:started:   inputs: " & " call72_994 = "& Convert_SLV_To_Hex_String(call72_994));
          --
        end if; 
        if type_cast_997_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_997_inst:finished:  outputs: " & " conv74_998= "  & Convert_SLV_To_Hex_String(conv74_998));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_997_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_997_inst_req_0;
      type_cast_997_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_997_inst_req_1;
      type_cast_997_inst_ack_1<= rack(0);
      type_cast_997_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_997_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call72_994,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_998,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_1221_index_1_rename flow-through 
    process(R_ix_x1x_xlcssa_1220_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_1221_index_1_rename:flowthrough  inputs: " & " R_ix_x1x_xlcssa_1220_resized = "& Convert_SLV_To_Hex_String(R_ix_x1x_xlcssa_1220_resized) & "outputs: " & " R_ix_x1x_xlcssa_1220_scaled= "  & Convert_SLV_To_Hex_String(R_ix_x1x_xlcssa_1220_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1221_index_1_rename
    process(R_ix_x1x_xlcssa_1220_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_1220_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_1220_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1221_index_1_resize flow-through 
    process(R_ix_x1x_xlcssa_1220_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_1221_index_1_resize:flowthrough  inputs: " & " ix_x1x_xlcssa_1086 = "& Convert_SLV_To_Hex_String(ix_x1x_xlcssa_1086) & "outputs: " & " R_ix_x1x_xlcssa_1220_resized= "  & Convert_SLV_To_Hex_String(R_ix_x1x_xlcssa_1220_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1221_index_1_resize
    process(ix_x1x_xlcssa_1086) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_1086;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_1220_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1221_root_address_inst flow-through 
    process(array_obj_ref_1221_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_1221_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1221_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1221_final_offset) & "outputs: " & " array_obj_ref_1221_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1221_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1221_root_address_inst
    process(array_obj_ref_1221_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1221_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1221_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_587_index_1_rename flow-through 
    process(R_indvar256_586_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_587_index_1_rename:flowthrough  inputs: " & " R_indvar256_586_resized = "& Convert_SLV_To_Hex_String(R_indvar256_586_resized) & "outputs: " & " R_indvar256_586_scaled= "  & Convert_SLV_To_Hex_String(R_indvar256_586_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_587_index_1_rename
    process(R_indvar256_586_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar256_586_resized;
      ov(13 downto 0) := iv;
      R_indvar256_586_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_587_index_1_resize flow-through 
    process(R_indvar256_586_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_587_index_1_resize:flowthrough  inputs: " & " indvar256_575 = "& Convert_SLV_To_Hex_String(indvar256_575) & "outputs: " & " R_indvar256_586_resized= "  & Convert_SLV_To_Hex_String(R_indvar256_586_resized));
      --
    end process; 
    -- equivalence array_obj_ref_587_index_1_resize
    process(indvar256_575) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar256_575;
      ov := iv(13 downto 0);
      R_indvar256_586_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_587_root_address_inst flow-through 
    process(array_obj_ref_587_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_587_root_address_inst:flowthrough  inputs: " & " array_obj_ref_587_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_587_final_offset) & "outputs: " & " array_obj_ref_587_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_587_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_587_root_address_inst
    process(array_obj_ref_587_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_587_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_587_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_827_index_1_rename flow-through 
    process(R_ix_x0x_xlcssa_826_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_827_index_1_rename:flowthrough  inputs: " & " R_ix_x0x_xlcssa_826_resized = "& Convert_SLV_To_Hex_String(R_ix_x0x_xlcssa_826_resized) & "outputs: " & " R_ix_x0x_xlcssa_826_scaled= "  & Convert_SLV_To_Hex_String(R_ix_x0x_xlcssa_826_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_827_index_1_rename
    process(R_ix_x0x_xlcssa_826_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_826_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_826_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_827_index_1_resize flow-through 
    process(R_ix_x0x_xlcssa_826_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_827_index_1_resize:flowthrough  inputs: " & " ix_x0x_xlcssa_697 = "& Convert_SLV_To_Hex_String(ix_x0x_xlcssa_697) & "outputs: " & " R_ix_x0x_xlcssa_826_resized= "  & Convert_SLV_To_Hex_String(R_ix_x0x_xlcssa_826_resized));
      --
    end process; 
    -- equivalence array_obj_ref_827_index_1_resize
    process(ix_x0x_xlcssa_697) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_697;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_826_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_827_root_address_inst flow-through 
    process(array_obj_ref_827_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_827_root_address_inst:flowthrough  inputs: " & " array_obj_ref_827_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_827_final_offset) & "outputs: " & " array_obj_ref_827_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_827_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_827_root_address_inst
    process(array_obj_ref_827_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_827_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_827_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_976_index_1_rename flow-through 
    process(R_indvar240_975_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_976_index_1_rename:flowthrough  inputs: " & " R_indvar240_975_resized = "& Convert_SLV_To_Hex_String(R_indvar240_975_resized) & "outputs: " & " R_indvar240_975_scaled= "  & Convert_SLV_To_Hex_String(R_indvar240_975_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_976_index_1_rename
    process(R_indvar240_975_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar240_975_resized;
      ov(13 downto 0) := iv;
      R_indvar240_975_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_976_index_1_resize flow-through 
    process(R_indvar240_975_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_976_index_1_resize:flowthrough  inputs: " & " indvar240_964 = "& Convert_SLV_To_Hex_String(indvar240_964) & "outputs: " & " R_indvar240_975_resized= "  & Convert_SLV_To_Hex_String(R_indvar240_975_resized));
      --
    end process; 
    -- equivalence array_obj_ref_976_index_1_resize
    process(indvar240_964) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar240_964;
      ov := iv(13 downto 0);
      R_indvar240_975_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_976_root_address_inst flow-through 
    process(array_obj_ref_976_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_976_root_address_inst:flowthrough  inputs: " & " array_obj_ref_976_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_976_final_offset) & "outputs: " & " array_obj_ref_976_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_976_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_976_root_address_inst
    process(array_obj_ref_976_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_976_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_976_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1041_addr_0 flow-through 
    process(ptr_deref_1041_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_1041_addr_0:flowthrough  inputs: " & " ptr_deref_1041_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1041_root_address) & "outputs: " & " ptr_deref_1041_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1041_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_1041_addr_0
    process(ptr_deref_1041_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1041_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1041_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1041_base_resize flow-through 
    process(ptr_deref_1041_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_1041_base_resize:flowthrough  inputs: " & " arrayidx91_978 = "& Convert_SLV_To_Hex_String(arrayidx91_978) & "outputs: " & " ptr_deref_1041_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1041_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_1041_base_resize
    process(arrayidx91_978) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx91_978;
      ov := iv(13 downto 0);
      ptr_deref_1041_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1041_gather_scatter flow-through 
    process(ptr_deref_1041_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_1041_gather_scatter:flowthrough  inputs: " & " add87_1039 = "& Convert_SLV_To_Hex_String(add87_1039) & "outputs: " & " ptr_deref_1041_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1041_data_0));
      --
    end process; 
    -- equivalence ptr_deref_1041_gather_scatter
    process(add87_1039) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add87_1039;
      ov(63 downto 0) := iv;
      ptr_deref_1041_data_0 <= ov(63 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1041_root_address_inst flow-through 
    process(ptr_deref_1041_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_1041_root_address_inst:flowthrough  inputs: " & " ptr_deref_1041_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_1041_resized_base_address) & "outputs: " & " ptr_deref_1041_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1041_root_address));
      --
    end process; 
    -- equivalence ptr_deref_1041_root_address_inst
    process(ptr_deref_1041_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1041_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1041_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1225_addr_0 flow-through 
    process(ptr_deref_1225_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_1225_addr_0:flowthrough  inputs: " & " ptr_deref_1225_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1225_root_address) & "outputs: " & " ptr_deref_1225_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1225_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_1225_addr_0
    process(ptr_deref_1225_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1225_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1225_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1225_base_resize flow-through 
    process(ptr_deref_1225_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_1225_base_resize:flowthrough  inputs: " & " arrayidx106_1223 = "& Convert_SLV_To_Hex_String(arrayidx106_1223) & "outputs: " & " ptr_deref_1225_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1225_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_1225_base_resize
    process(arrayidx106_1223) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx106_1223;
      ov := iv(13 downto 0);
      ptr_deref_1225_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1225_gather_scatter flow-through 
    process(ptr_deref_1225_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_1225_gather_scatter:flowthrough  inputs: " & " shl12x_xi187_1216 = "& Convert_SLV_To_Hex_String(shl12x_xi187_1216) & "outputs: " & " ptr_deref_1225_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1225_data_0));
      --
    end process; 
    -- equivalence ptr_deref_1225_gather_scatter
    process(shl12x_xi187_1216) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl12x_xi187_1216;
      ov(63 downto 0) := iv;
      ptr_deref_1225_data_0 <= ov(63 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1225_root_address_inst flow-through 
    process(ptr_deref_1225_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_1225_root_address_inst:flowthrough  inputs: " & " ptr_deref_1225_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_1225_resized_base_address) & "outputs: " & " ptr_deref_1225_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1225_root_address));
      --
    end process; 
    -- equivalence ptr_deref_1225_root_address_inst
    process(ptr_deref_1225_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1225_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1225_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_652_addr_0 flow-through 
    process(ptr_deref_652_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_652_addr_0:flowthrough  inputs: " & " ptr_deref_652_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_652_root_address) & "outputs: " & " ptr_deref_652_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_652_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_652_addr_0
    process(ptr_deref_652_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_652_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_652_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_652_base_resize flow-through 
    process(ptr_deref_652_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_652_base_resize:flowthrough  inputs: " & " arrayidx_589 = "& Convert_SLV_To_Hex_String(arrayidx_589) & "outputs: " & " ptr_deref_652_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_652_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_652_base_resize
    process(arrayidx_589) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_589;
      ov := iv(13 downto 0);
      ptr_deref_652_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_652_gather_scatter flow-through 
    process(ptr_deref_652_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_652_gather_scatter:flowthrough  inputs: " & " add36_650 = "& Convert_SLV_To_Hex_String(add36_650) & "outputs: " & " ptr_deref_652_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_652_data_0));
      --
    end process; 
    -- equivalence ptr_deref_652_gather_scatter
    process(add36_650) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add36_650;
      ov(63 downto 0) := iv;
      ptr_deref_652_data_0 <= ov(63 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_652_root_address_inst flow-through 
    process(ptr_deref_652_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_652_root_address_inst:flowthrough  inputs: " & " ptr_deref_652_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_652_resized_base_address) & "outputs: " & " ptr_deref_652_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_652_root_address));
      --
    end process; 
    -- equivalence ptr_deref_652_root_address_inst
    process(ptr_deref_652_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_652_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_652_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_831_addr_0 flow-through 
    process(ptr_deref_831_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_831_addr_0:flowthrough  inputs: " & " ptr_deref_831_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_831_root_address) & "outputs: " & " ptr_deref_831_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_831_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_831_addr_0
    process(ptr_deref_831_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_831_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_831_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_831_base_resize flow-through 
    process(ptr_deref_831_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_831_base_resize:flowthrough  inputs: " & " arrayidx47_829 = "& Convert_SLV_To_Hex_String(arrayidx47_829) & "outputs: " & " ptr_deref_831_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_831_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_831_base_resize
    process(arrayidx47_829) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx47_829;
      ov := iv(13 downto 0);
      ptr_deref_831_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_831_gather_scatter flow-through 
    process(ptr_deref_831_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_831_gather_scatter:flowthrough  inputs: " & " shl12x_xi_822 = "& Convert_SLV_To_Hex_String(shl12x_xi_822) & "outputs: " & " ptr_deref_831_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_831_data_0));
      --
    end process; 
    -- equivalence ptr_deref_831_gather_scatter
    process(shl12x_xi_822) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl12x_xi_822;
      ov(63 downto 0) := iv;
      ptr_deref_831_data_0 <= ov(63 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_831_root_address_inst flow-through 
    process(ptr_deref_831_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_831_root_address_inst:flowthrough  inputs: " & " ptr_deref_831_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_831_resized_base_address) & "outputs: " & " ptr_deref_831_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_831_root_address));
      --
    end process; 
    -- equivalence ptr_deref_831_root_address_inst
    process(ptr_deref_831_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_831_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_831_root_address <= ov(13 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1055_branch_req_0," req0 if_stmt_1055_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1055_branch_ack_0," ack0 if_stmt_1055_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1055_branch_ack_1," ack1 if_stmt_1055_branch");
    if_stmt_1055_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond26_1054;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1055_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1055_branch_req_0,
          ack0 => if_stmt_1055_branch_ack_0,
          ack1 => if_stmt_1055_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1106_branch_req_0," req0 if_stmt_1106_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1106_branch_ack_0," ack0 if_stmt_1106_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1106_branch_ack_1," ack1 if_stmt_1106_branch");
    if_stmt_1106_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool98_1105;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1106_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1106_branch_req_0,
          ack0 => if_stmt_1106_branch_ack_0,
          ack1 => if_stmt_1106_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1182_branch_req_0," req0 if_stmt_1182_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1182_branch_ack_0," ack0 if_stmt_1182_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1182_branch_ack_1," ack1 if_stmt_1182_branch");
    if_stmt_1182_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1181;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1182_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1182_branch_req_0,
          ack0 => if_stmt_1182_branch_ack_0,
          ack1 => if_stmt_1182_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1346_branch_req_0," req0 if_stmt_1346_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1346_branch_ack_0," ack0 if_stmt_1346_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1346_branch_ack_1," ack1 if_stmt_1346_branch");
    if_stmt_1346_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond7_1345;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1346_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1346_branch_req_0,
          ack0 => if_stmt_1346_branch_ack_0,
          ack1 => if_stmt_1346_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_504_branch_req_0," req0 if_stmt_504_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_504_branch_ack_0," ack0 if_stmt_504_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_504_branch_ack_1," ack1 if_stmt_504_branch");
    if_stmt_504_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp195_503;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_504_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_504_branch_req_0,
          ack0 => if_stmt_504_branch_ack_0,
          ack1 => if_stmt_504_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_666_branch_req_0," req0 if_stmt_666_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_666_branch_ack_0," ack0 if_stmt_666_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_666_branch_ack_1," ack1 if_stmt_666_branch");
    if_stmt_666_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond37_665;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_666_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_666_branch_req_0,
          ack0 => if_stmt_666_branch_ack_0,
          ack1 => if_stmt_666_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_717_branch_req_0," req0 if_stmt_717_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_717_branch_ack_0," ack0 if_stmt_717_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_717_branch_ack_1," ack1 if_stmt_717_branch");
    if_stmt_717_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_716;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_717_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_717_branch_req_0,
          ack0 => if_stmt_717_branch_ack_0,
          ack1 => if_stmt_717_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_788_branch_req_0," req0 if_stmt_788_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_788_branch_ack_0," ack0 if_stmt_788_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_788_branch_ack_1," ack1 if_stmt_788_branch");
    if_stmt_788_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_787;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_788_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_788_branch_req_0,
          ack0 => if_stmt_788_branch_ack_0,
          ack1 => if_stmt_788_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_884_branch_req_0," req0 if_stmt_884_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_884_branch_ack_0," ack0 if_stmt_884_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_884_branch_ack_1," ack1 if_stmt_884_branch");
    if_stmt_884_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp65191_883;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_884_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_884_branch_req_0,
          ack0 => if_stmt_884_branch_ack_0,
          ack1 => if_stmt_884_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u16_u16_1175_inst flow-through 
    process(incx_xi179_1176) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ADD_u16_u16_1175_inst:flowthrough inputs: " & " nx_x016x_xi173_1138 = "& Convert_SLV_To_Hex_String(nx_x016x_xi173_1138) & " type_cast_1174_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1174_wire_constant) & " outputs:" & " incx_xi179_1176= "  & Convert_SLV_To_Hex_String(incx_xi179_1176));
      --
    end process; 
    -- binary operator ADD_u16_u16_1175_inst
    process(nx_x016x_xi173_1138) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x016x_xi173_1138, type_cast_1174_wire_constant, tmp_var);
      incx_xi179_1176 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1255_inst flow-through 
    process(sub_1256) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ADD_u16_u16_1255_inst:flowthrough inputs: " & " call4_450 = "& Convert_SLV_To_Hex_String(call4_450) & " type_cast_1254_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1254_wire_constant) & " outputs:" & " sub_1256= "  & Convert_SLV_To_Hex_String(sub_1256));
      --
    end process; 
    -- binary operator ADD_u16_u16_1255_inst
    process(call4_450) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call4_450, type_cast_1254_wire_constant, tmp_var);
      sub_1256 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1261_inst flow-through 
    process(sub149_1262) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ADD_u16_u16_1261_inst:flowthrough inputs: " & " call6_456 = "& Convert_SLV_To_Hex_String(call6_456) & " type_cast_1260_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1260_wire_constant) & " outputs:" & " sub149_1262= "  & Convert_SLV_To_Hex_String(sub149_1262));
      --
    end process; 
    -- binary operator ADD_u16_u16_1261_inst
    process(call6_456) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call6_456, type_cast_1260_wire_constant, tmp_var);
      sub149_1262 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1267_inst flow-through 
    process(tmp216_1268) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ADD_u16_u16_1267_inst:flowthrough inputs: " & " call5_453 = "& Convert_SLV_To_Hex_String(call5_453) & " type_cast_1266_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1266_wire_constant) & " outputs:" & " tmp216_1268= "  & Convert_SLV_To_Hex_String(tmp216_1268));
      --
    end process; 
    -- binary operator ADD_u16_u16_1267_inst
    process(call5_453) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call5_453, type_cast_1266_wire_constant, tmp_var);
      tmp216_1268 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_781_inst flow-through 
    process(incx_xi_782) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ADD_u16_u16_781_inst:flowthrough inputs: " & " nx_x016x_xi_744 = "& Convert_SLV_To_Hex_String(nx_x016x_xi_744) & " type_cast_780_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_780_wire_constant) & " outputs:" & " incx_xi_782= "  & Convert_SLV_To_Hex_String(incx_xi_782));
      --
    end process; 
    -- binary operator ADD_u16_u16_781_inst
    process(nx_x016x_xi_744) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x016x_xi_744, type_cast_780_wire_constant, tmp_var);
      incx_xi_782 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1277_inst flow-through 
    process(tmp6_1278) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ADD_u32_u32_1277_inst:flowthrough inputs: " & " tmp5_1272 = "& Convert_SLV_To_Hex_String(tmp5_1272) & " type_cast_1276_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1276_wire_constant) & " outputs:" & " tmp6_1278= "  & Convert_SLV_To_Hex_String(tmp6_1278));
      --
    end process; 
    -- binary operator ADD_u32_u32_1277_inst
    process(tmp5_1272) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_1272, type_cast_1276_wire_constant, tmp_var);
      tmp6_1278 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1315_inst flow-through 
    process(mul140_1316) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ADD_u32_u32_1315_inst:flowthrough inputs: " & " tmp11_1296 = "& Convert_SLV_To_Hex_String(tmp11_1296) & " mul134_1311 = "& Convert_SLV_To_Hex_String(mul134_1311) & " outputs:" & " mul140_1316= "  & Convert_SLV_To_Hex_String(mul140_1316));
      --
    end process; 
    -- binary operator ADD_u32_u32_1315_inst
    process(tmp11_1296, mul134_1311) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp11_1296, mul134_1311, tmp_var);
      mul140_1316 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1339_inst flow-through 
    process(indvarx_xnext_1340) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ADD_u32_u32_1339_inst:flowthrough inputs: " & " indvar_1299 = "& Convert_SLV_To_Hex_String(indvar_1299) & " type_cast_1338_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1338_wire_constant) & " outputs:" & " indvarx_xnext_1340= "  & Convert_SLV_To_Hex_String(indvarx_xnext_1340));
      --
    end process; 
    -- binary operator ADD_u32_u32_1339_inst
    process(indvar_1299) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1299, type_cast_1338_wire_constant, tmp_var);
      indvarx_xnext_1340 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u64_u64_1048_inst flow-through 
    process(indvarx_xnext241_1049) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ADD_u64_u64_1048_inst:flowthrough inputs: " & " indvar240_964 = "& Convert_SLV_To_Hex_String(indvar240_964) & " type_cast_1047_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1047_wire_constant) & " outputs:" & " indvarx_xnext241_1049= "  & Convert_SLV_To_Hex_String(indvarx_xnext241_1049));
      --
    end process; 
    -- binary operator ADD_u64_u64_1048_inst
    process(indvar240_964) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar240_964, type_cast_1047_wire_constant, tmp_var);
      indvarx_xnext241_1049 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u64_u64_659_inst flow-through 
    process(indvarx_xnext257_660) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ADD_u64_u64_659_inst:flowthrough inputs: " & " indvar256_575 = "& Convert_SLV_To_Hex_String(indvar256_575) & " type_cast_658_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_658_wire_constant) & " outputs:" & " indvarx_xnext257_660= "  & Convert_SLV_To_Hex_String(indvarx_xnext257_660));
      --
    end process; 
    -- binary operator ADD_u64_u64_659_inst
    process(indvar256_575) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar256_575, type_cast_658_wire_constant, tmp_var);
      indvarx_xnext257_660 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u64_u64_1098_inst flow-through 
    process(and97_1099) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:AND_u64_u64_1098_inst:flowthrough inputs: " & " conv59_877 = "& Convert_SLV_To_Hex_String(conv59_877) & " type_cast_1097_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1097_wire_constant) & " outputs:" & " and97_1099= "  & Convert_SLV_To_Hex_String(and97_1099));
      --
    end process; 
    -- binary operator AND_u64_u64_1098_inst
    process(conv59_877) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv59_877, type_cast_1097_wire_constant, tmp_var);
      and97_1099 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u64_u64_1204_inst flow-through 
    process(mulx_xi185_1205) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:AND_u64_u64_1204_inst:flowthrough inputs: " & " iNsTr_52_1199 = "& Convert_SLV_To_Hex_String(iNsTr_52_1199) & " type_cast_1203_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1203_wire_constant) & " outputs:" & " mulx_xi185_1205= "  & Convert_SLV_To_Hex_String(mulx_xi185_1205));
      --
    end process; 
    -- binary operator AND_u64_u64_1204_inst
    process(iNsTr_52_1199) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_52_1199, type_cast_1203_wire_constant, tmp_var);
      mulx_xi185_1205 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u64_u64_709_inst flow-through 
    process(and_710) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:AND_u64_u64_709_inst:flowthrough inputs: " & " conv13_497 = "& Convert_SLV_To_Hex_String(conv13_497) & " type_cast_708_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_708_wire_constant) & " outputs:" & " and_710= "  & Convert_SLV_To_Hex_String(and_710));
      --
    end process; 
    -- binary operator AND_u64_u64_709_inst
    process(conv13_497) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv13_497, type_cast_708_wire_constant, tmp_var);
      and_710 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u64_u64_810_inst flow-through 
    process(mulx_xi_811) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:AND_u64_u64_810_inst:flowthrough inputs: " & " iNsTr_38_805 = "& Convert_SLV_To_Hex_String(iNsTr_38_805) & " type_cast_809_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_809_wire_constant) & " outputs:" & " mulx_xi_811= "  & Convert_SLV_To_Hex_String(mulx_xi_811));
      --
    end process; 
    -- binary operator AND_u64_u64_810_inst
    process(iNsTr_38_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_38_805, type_cast_809_wire_constant, tmp_var);
      mulx_xi_811 <= tmp_var; --
    end process;
    -- logger for split-operator ASHR_i64_i64_1081_inst flow-through 
    process(ASHR_i64_i64_1081_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ASHR_i64_i64_1081_inst:flowthrough inputs: " & " type_cast_1077_wire = "& Convert_SLV_To_Hex_String(type_cast_1077_wire) & " type_cast_1080_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1080_wire_constant) & " outputs:" & " ASHR_i64_i64_1081_wire= "  & Convert_SLV_To_Hex_String(ASHR_i64_i64_1081_wire));
      --
    end process; 
    -- binary operator ASHR_i64_i64_1081_inst
    process(type_cast_1077_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1077_wire, type_cast_1080_wire_constant, tmp_var);
      ASHR_i64_i64_1081_wire <= tmp_var; --
    end process;
    -- logger for split-operator ASHR_i64_i64_495_inst flow-through 
    process(ASHR_i64_i64_495_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ASHR_i64_i64_495_inst:flowthrough inputs: " & " type_cast_491_wire = "& Convert_SLV_To_Hex_String(type_cast_491_wire) & " type_cast_494_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_494_wire_constant) & " outputs:" & " ASHR_i64_i64_495_wire= "  & Convert_SLV_To_Hex_String(ASHR_i64_i64_495_wire));
      --
    end process; 
    -- binary operator ASHR_i64_i64_495_inst
    process(type_cast_491_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_491_wire, type_cast_494_wire_constant, tmp_var);
      ASHR_i64_i64_495_wire <= tmp_var; --
    end process;
    -- logger for split-operator ASHR_i64_i64_692_inst flow-through 
    process(ASHR_i64_i64_692_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ASHR_i64_i64_692_inst:flowthrough inputs: " & " type_cast_688_wire = "& Convert_SLV_To_Hex_String(type_cast_688_wire) & " type_cast_691_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_691_wire_constant) & " outputs:" & " ASHR_i64_i64_692_wire= "  & Convert_SLV_To_Hex_String(ASHR_i64_i64_692_wire));
      --
    end process; 
    -- binary operator ASHR_i64_i64_692_inst
    process(type_cast_688_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_688_wire, type_cast_691_wire_constant, tmp_var);
      ASHR_i64_i64_692_wire <= tmp_var; --
    end process;
    -- logger for split-operator ASHR_i64_i64_875_inst flow-through 
    process(ASHR_i64_i64_875_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ASHR_i64_i64_875_inst:flowthrough inputs: " & " type_cast_871_wire = "& Convert_SLV_To_Hex_String(type_cast_871_wire) & " type_cast_874_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_874_wire_constant) & " outputs:" & " ASHR_i64_i64_875_wire= "  & Convert_SLV_To_Hex_String(ASHR_i64_i64_875_wire));
      --
    end process; 
    -- binary operator ASHR_i64_i64_875_inst
    process(type_cast_871_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_871_wire, type_cast_874_wire_constant, tmp_var);
      ASHR_i64_i64_875_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u16_u1_1180_inst flow-through 
    process(exitcond_1181) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:EQ_u16_u1_1180_inst:flowthrough inputs: " & " incx_xi179_1176 = "& Convert_SLV_To_Hex_String(incx_xi179_1176) & " tmp4_1135 = "& Convert_SLV_To_Hex_String(tmp4_1135) & " outputs:" & " exitcond_1181= "  & Convert_SLV_To_Hex_String(exitcond_1181));
      --
    end process; 
    -- binary operator EQ_u16_u1_1180_inst
    process(incx_xi179_1176, tmp4_1135) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(incx_xi179_1176, tmp4_1135, tmp_var);
      exitcond_1181 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u16_u1_786_inst flow-through 
    process(exitcond2_787) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:EQ_u16_u1_786_inst:flowthrough inputs: " & " incx_xi_782 = "& Convert_SLV_To_Hex_String(incx_xi_782) & " tmp1_741 = "& Convert_SLV_To_Hex_String(tmp1_741) & " outputs:" & " exitcond2_787= "  & Convert_SLV_To_Hex_String(exitcond2_787));
      --
    end process; 
    -- binary operator EQ_u16_u1_786_inst
    process(incx_xi_782, tmp1_741) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(incx_xi_782, tmp1_741, tmp_var);
      exitcond2_787 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u32_u1_1344_inst flow-through 
    process(exitcond7_1345) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:EQ_u32_u1_1344_inst:flowthrough inputs: " & " indvarx_xnext_1340 = "& Convert_SLV_To_Hex_String(indvarx_xnext_1340) & " tmp6_1278 = "& Convert_SLV_To_Hex_String(tmp6_1278) & " outputs:" & " exitcond7_1345= "  & Convert_SLV_To_Hex_String(exitcond7_1345));
      --
    end process; 
    -- binary operator EQ_u32_u1_1344_inst
    process(indvarx_xnext_1340, tmp6_1278) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1340, tmp6_1278, tmp_var);
      exitcond7_1345 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u64_u1_1053_inst flow-through 
    process(exitcond26_1054) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:EQ_u64_u1_1053_inst:flowthrough inputs: " & " indvarx_xnext241_1049 = "& Convert_SLV_To_Hex_String(indvarx_xnext241_1049) & " umax25_961 = "& Convert_SLV_To_Hex_String(umax25_961) & " outputs:" & " exitcond26_1054= "  & Convert_SLV_To_Hex_String(exitcond26_1054));
      --
    end process; 
    -- binary operator EQ_u64_u1_1053_inst
    process(indvarx_xnext241_1049, umax25_961) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext241_1049, umax25_961, tmp_var);
      exitcond26_1054 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u64_u1_1104_inst flow-through 
    process(tobool98_1105) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:EQ_u64_u1_1104_inst:flowthrough inputs: " & " and97_1099 = "& Convert_SLV_To_Hex_String(and97_1099) & " type_cast_1103_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1103_wire_constant) & " outputs:" & " tobool98_1105= "  & Convert_SLV_To_Hex_String(tobool98_1105));
      --
    end process; 
    -- binary operator EQ_u64_u1_1104_inst
    process(and97_1099) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and97_1099, type_cast_1103_wire_constant, tmp_var);
      tobool98_1105 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u64_u1_664_inst flow-through 
    process(exitcond37_665) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:EQ_u64_u1_664_inst:flowthrough inputs: " & " indvarx_xnext257_660 = "& Convert_SLV_To_Hex_String(indvarx_xnext257_660) & " umax36_572 = "& Convert_SLV_To_Hex_String(umax36_572) & " outputs:" & " exitcond37_665= "  & Convert_SLV_To_Hex_String(exitcond37_665));
      --
    end process; 
    -- binary operator EQ_u64_u1_664_inst
    process(indvarx_xnext257_660, umax36_572) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext257_660, umax36_572, tmp_var);
      exitcond37_665 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u64_u1_715_inst flow-through 
    process(tobool_716) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:EQ_u64_u1_715_inst:flowthrough inputs: " & " and_710 = "& Convert_SLV_To_Hex_String(and_710) & " type_cast_714_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_714_wire_constant) & " outputs:" & " tobool_716= "  & Convert_SLV_To_Hex_String(tobool_716));
      --
    end process; 
    -- binary operator EQ_u64_u1_715_inst
    process(and_710) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_710, type_cast_714_wire_constant, tmp_var);
      tobool_716 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u64_u64_515_inst flow-through 
    process(tmp250_516) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:LSHR_u64_u64_515_inst:flowthrough inputs: " & " conv13_497 = "& Convert_SLV_To_Hex_String(conv13_497) & " type_cast_514_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_514_wire_constant) & " outputs:" & " tmp250_516= "  & Convert_SLV_To_Hex_String(tmp250_516));
      --
    end process; 
    -- binary operator LSHR_u64_u64_515_inst
    process(conv13_497) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv13_497, type_cast_514_wire_constant, tmp_var);
      tmp250_516 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u64_u64_558_inst flow-through 
    process(tmp34_559) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:LSHR_u64_u64_558_inst:flowthrough inputs: " & " tmp33_553 = "& Convert_SLV_To_Hex_String(tmp33_553) & " type_cast_557_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_557_wire_constant) & " outputs:" & " tmp34_559= "  & Convert_SLV_To_Hex_String(tmp34_559));
      --
    end process; 
    -- binary operator LSHR_u64_u64_558_inst
    process(tmp33_553) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp33_553, type_cast_557_wire_constant, tmp_var);
      tmp34_559 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u64_u64_895_inst flow-through 
    process(tmp235_896) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:LSHR_u64_u64_895_inst:flowthrough inputs: " & " conv59_877 = "& Convert_SLV_To_Hex_String(conv59_877) & " type_cast_894_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_894_wire_constant) & " outputs:" & " tmp235_896= "  & Convert_SLV_To_Hex_String(tmp235_896));
      --
    end process; 
    -- binary operator LSHR_u64_u64_895_inst
    process(conv59_877) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv59_877, type_cast_894_wire_constant, tmp_var);
      tmp235_896 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u64_u64_947_inst flow-through 
    process(tmp23_948) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:LSHR_u64_u64_947_inst:flowthrough inputs: " & " tmp22_942 = "& Convert_SLV_To_Hex_String(tmp22_942) & " type_cast_946_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_946_wire_constant) & " outputs:" & " tmp23_948= "  & Convert_SLV_To_Hex_String(tmp23_948));
      --
    end process; 
    -- binary operator LSHR_u64_u64_947_inst
    process(tmp22_942) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp22_942, type_cast_946_wire_constant, tmp_var);
      tmp23_948 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1116_inst flow-through 
    process(tmp208_1117) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u16_u16_1116_inst:flowthrough inputs: " & " call5_453 = "& Convert_SLV_To_Hex_String(call5_453) & " call2_444 = "& Convert_SLV_To_Hex_String(call2_444) & " outputs:" & " tmp208_1117= "  & Convert_SLV_To_Hex_String(tmp208_1117));
      --
    end process; 
    -- binary operator MUL_u16_u16_1116_inst
    process(call5_453, call2_444) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call5_453, call2_444, tmp_var);
      tmp208_1117 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1121_inst flow-through 
    process(tmp210_1122) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u16_u16_1121_inst:flowthrough inputs: " & " tmp208_1117 = "& Convert_SLV_To_Hex_String(tmp208_1117) & " call6_456 = "& Convert_SLV_To_Hex_String(call6_456) & " outputs:" & " tmp210_1122= "  & Convert_SLV_To_Hex_String(tmp210_1122));
      --
    end process; 
    -- binary operator MUL_u16_u16_1121_inst
    process(tmp208_1117, call6_456) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp208_1117, call6_456, tmp_var);
      tmp210_1122 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1126_inst flow-through 
    process(tmp212_1127) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u16_u16_1126_inst:flowthrough inputs: " & " tmp210_1122 = "& Convert_SLV_To_Hex_String(tmp210_1122) & " call7_459 = "& Convert_SLV_To_Hex_String(call7_459) & " outputs:" & " tmp212_1127= "  & Convert_SLV_To_Hex_String(tmp212_1127));
      --
    end process; 
    -- binary operator MUL_u16_u16_1126_inst
    process(tmp210_1122, call7_459) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp210_1122, call7_459, tmp_var);
      tmp212_1127 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1237_inst flow-through 
    process(mul116_1238) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u16_u16_1237_inst:flowthrough inputs: " & " call7_459 = "& Convert_SLV_To_Hex_String(call7_459) & " call2_444 = "& Convert_SLV_To_Hex_String(call2_444) & " outputs:" & " mul116_1238= "  & Convert_SLV_To_Hex_String(mul116_1238));
      --
    end process; 
    -- binary operator MUL_u16_u16_1237_inst
    process(call7_459, call2_444) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call7_459, call2_444, tmp_var);
      mul116_1238 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1242_inst flow-through 
    process(mul129_1243) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u16_u16_1242_inst:flowthrough inputs: " & " call4_450 = "& Convert_SLV_To_Hex_String(call4_450) & " call3_447 = "& Convert_SLV_To_Hex_String(call3_447) & " outputs:" & " mul129_1243= "  & Convert_SLV_To_Hex_String(mul129_1243));
      --
    end process; 
    -- binary operator MUL_u16_u16_1242_inst
    process(call4_450, call3_447) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call4_450, call3_447, tmp_var);
      mul129_1243 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1286_inst flow-through 
    process(tmp9_1287) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u16_u16_1286_inst:flowthrough inputs: " & " call7_459 = "& Convert_SLV_To_Hex_String(call7_459) & " call2_444 = "& Convert_SLV_To_Hex_String(call2_444) & " outputs:" & " tmp9_1287= "  & Convert_SLV_To_Hex_String(tmp9_1287));
      --
    end process; 
    -- binary operator MUL_u16_u16_1286_inst
    process(call7_459, call2_444) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call7_459, call2_444, tmp_var);
      tmp9_1287 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_727_inst flow-through 
    process(tmp201_728) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u16_u16_727_inst:flowthrough inputs: " & " call1_441 = "& Convert_SLV_To_Hex_String(call1_441) & " call_438 = "& Convert_SLV_To_Hex_String(call_438) & " outputs:" & " tmp201_728= "  & Convert_SLV_To_Hex_String(tmp201_728));
      --
    end process; 
    -- binary operator MUL_u16_u16_727_inst
    process(call1_441, call_438) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call1_441, call_438, tmp_var);
      tmp201_728 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_732_inst flow-through 
    process(tmp203_733) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u16_u16_732_inst:flowthrough inputs: " & " tmp201_728 = "& Convert_SLV_To_Hex_String(tmp201_728) & " call2_444 = "& Convert_SLV_To_Hex_String(call2_444) & " outputs:" & " tmp203_733= "  & Convert_SLV_To_Hex_String(tmp203_733));
      --
    end process; 
    -- binary operator MUL_u16_u16_732_inst
    process(tmp201_728, call2_444) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp201_728, call2_444, tmp_var);
      tmp203_733 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u32_u32_1295_inst flow-through 
    process(tmp11_1296) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u32_u32_1295_inst:flowthrough inputs: " & " tmp8_1282 = "& Convert_SLV_To_Hex_String(tmp8_1282) & " tmp10_1291 = "& Convert_SLV_To_Hex_String(tmp10_1291) & " outputs:" & " tmp11_1296= "  & Convert_SLV_To_Hex_String(tmp11_1296));
      --
    end process; 
    -- binary operator MUL_u32_u32_1295_inst
    process(tmp8_1282, tmp10_1291) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp8_1282, tmp10_1291, tmp_var);
      tmp11_1296 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u32_u32_1310_inst flow-through 
    process(mul134_1311) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u32_u32_1310_inst:flowthrough inputs: " & " tmp11_1296 = "& Convert_SLV_To_Hex_String(tmp11_1296) & " indvar_1299 = "& Convert_SLV_To_Hex_String(indvar_1299) & " outputs:" & " mul134_1311= "  & Convert_SLV_To_Hex_String(mul134_1311));
      --
    end process; 
    -- binary operator MUL_u32_u32_1310_inst
    process(tmp11_1296, indvar_1299) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp11_1296, indvar_1299, tmp_var);
      mul134_1311 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u64_u64_475_inst flow-through 
    process(mul_476) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u64_u64_475_inst:flowthrough inputs: " & " conv9_467 = "& Convert_SLV_To_Hex_String(conv9_467) & " conv_463 = "& Convert_SLV_To_Hex_String(conv_463) & " outputs:" & " mul_476= "  & Convert_SLV_To_Hex_String(mul_476));
      --
    end process; 
    -- binary operator MUL_u64_u64_475_inst
    process(conv9_467, conv_463) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv9_467, conv_463, tmp_var);
      mul_476 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u64_u64_480_inst flow-through 
    process(mul12_481) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u64_u64_480_inst:flowthrough inputs: " & " mul_476 = "& Convert_SLV_To_Hex_String(mul_476) & " conv11_471 = "& Convert_SLV_To_Hex_String(conv11_471) & " outputs:" & " mul12_481= "  & Convert_SLV_To_Hex_String(mul12_481));
      --
    end process; 
    -- binary operator MUL_u64_u64_480_inst
    process(mul_476, conv11_471) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_476, conv11_471, tmp_var);
      mul12_481 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u64_u64_534_inst flow-through 
    process(tmp29_535) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u64_u64_534_inst:flowthrough inputs: " & " tmp27_526 = "& Convert_SLV_To_Hex_String(tmp27_526) & " tmp28_530 = "& Convert_SLV_To_Hex_String(tmp28_530) & " outputs:" & " tmp29_535= "  & Convert_SLV_To_Hex_String(tmp29_535));
      --
    end process; 
    -- binary operator MUL_u64_u64_534_inst
    process(tmp27_526, tmp28_530) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp27_526, tmp28_530, tmp_var);
      tmp29_535 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u64_u64_543_inst flow-through 
    process(tmp31_544) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u64_u64_543_inst:flowthrough inputs: " & " tmp29_535 = "& Convert_SLV_To_Hex_String(tmp29_535) & " tmp30_539 = "& Convert_SLV_To_Hex_String(tmp30_539) & " outputs:" & " tmp31_544= "  & Convert_SLV_To_Hex_String(tmp31_544));
      --
    end process; 
    -- binary operator MUL_u64_u64_543_inst
    process(tmp29_535, tmp30_539) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp29_535, tmp30_539, tmp_var);
      tmp31_544 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u64_u64_851_inst flow-through 
    process(mul52_852) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u64_u64_851_inst:flowthrough inputs: " & " conv57_847 = "& Convert_SLV_To_Hex_String(conv57_847) & " conv11_471 = "& Convert_SLV_To_Hex_String(conv11_471) & " outputs:" & " mul52_852= "  & Convert_SLV_To_Hex_String(mul52_852));
      --
    end process; 
    -- binary operator MUL_u64_u64_851_inst
    process(conv57_847, conv11_471) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv57_847, conv11_471, tmp_var);
      mul52_852 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u64_u64_856_inst flow-through 
    process(mul55_857) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u64_u64_856_inst:flowthrough inputs: " & " mul52_852 = "& Convert_SLV_To_Hex_String(mul52_852) & " conv54_843 = "& Convert_SLV_To_Hex_String(conv54_843) & " outputs:" & " mul55_857= "  & Convert_SLV_To_Hex_String(mul55_857));
      --
    end process; 
    -- binary operator MUL_u64_u64_856_inst
    process(mul52_852, conv54_843) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul52_852, conv54_843, tmp_var);
      mul55_857 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u64_u64_861_inst flow-through 
    process(mul58_862) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u64_u64_861_inst:flowthrough inputs: " & " mul55_857 = "& Convert_SLV_To_Hex_String(mul55_857) & " conv51_839 = "& Convert_SLV_To_Hex_String(conv51_839) & " outputs:" & " mul58_862= "  & Convert_SLV_To_Hex_String(mul58_862));
      --
    end process; 
    -- binary operator MUL_u64_u64_861_inst
    process(mul55_857, conv51_839) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul55_857, conv51_839, tmp_var);
      mul58_862 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u64_u64_914_inst flow-through 
    process(tmp16_915) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u64_u64_914_inst:flowthrough inputs: " & " tmp14_906 = "& Convert_SLV_To_Hex_String(tmp14_906) & " tmp15_910 = "& Convert_SLV_To_Hex_String(tmp15_910) & " outputs:" & " tmp16_915= "  & Convert_SLV_To_Hex_String(tmp16_915));
      --
    end process; 
    -- binary operator MUL_u64_u64_914_inst
    process(tmp14_906, tmp15_910) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_906, tmp15_910, tmp_var);
      tmp16_915 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u64_u64_923_inst flow-through 
    process(tmp18_924) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u64_u64_923_inst:flowthrough inputs: " & " tmp16_915 = "& Convert_SLV_To_Hex_String(tmp16_915) & " tmp17_919 = "& Convert_SLV_To_Hex_String(tmp17_919) & " outputs:" & " tmp18_924= "  & Convert_SLV_To_Hex_String(tmp18_924));
      --
    end process; 
    -- binary operator MUL_u64_u64_923_inst
    process(tmp16_915, tmp17_919) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_915, tmp17_919, tmp_var);
      tmp18_924 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u64_u64_932_inst flow-through 
    process(tmp20_933) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:MUL_u64_u64_932_inst:flowthrough inputs: " & " tmp18_924 = "& Convert_SLV_To_Hex_String(tmp18_924) & " tmp19_928 = "& Convert_SLV_To_Hex_String(tmp19_928) & " outputs:" & " tmp20_933= "  & Convert_SLV_To_Hex_String(tmp20_933));
      --
    end process; 
    -- binary operator MUL_u64_u64_932_inst
    process(tmp18_924, tmp19_928) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp18_924, tmp19_928, tmp_var);
      tmp20_933 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u64_u64_1002_inst flow-through 
    process(add75_1003) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:OR_u64_u64_1002_inst:flowthrough inputs: " & " shl71_991 = "& Convert_SLV_To_Hex_String(shl71_991) & " conv74_998 = "& Convert_SLV_To_Hex_String(conv74_998) & " outputs:" & " add75_1003= "  & Convert_SLV_To_Hex_String(add75_1003));
      --
    end process; 
    -- binary operator OR_u64_u64_1002_inst
    process(shl71_991, conv74_998) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl71_991, conv74_998, tmp_var);
      add75_1003 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u64_u64_1020_inst flow-through 
    process(add81_1021) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:OR_u64_u64_1020_inst:flowthrough inputs: " & " shl77_1009 = "& Convert_SLV_To_Hex_String(shl77_1009) & " conv80_1016 = "& Convert_SLV_To_Hex_String(conv80_1016) & " outputs:" & " add81_1021= "  & Convert_SLV_To_Hex_String(add81_1021));
      --
    end process; 
    -- binary operator OR_u64_u64_1020_inst
    process(shl77_1009, conv80_1016) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl77_1009, conv80_1016, tmp_var);
      add81_1021 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u64_u64_1038_inst flow-through 
    process(add87_1039) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:OR_u64_u64_1038_inst:flowthrough inputs: " & " shl83_1027 = "& Convert_SLV_To_Hex_String(shl83_1027) & " conv86_1034 = "& Convert_SLV_To_Hex_String(conv86_1034) & " outputs:" & " add87_1039= "  & Convert_SLV_To_Hex_String(add87_1039));
      --
    end process; 
    -- binary operator OR_u64_u64_1038_inst
    process(shl83_1027, conv86_1034) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl83_1027, conv86_1034, tmp_var);
      add87_1039 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u64_u64_1163_inst flow-through 
    process(addx_xi177_1164) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:OR_u64_u64_1163_inst:flowthrough inputs: " & " conv5x_xi176_1159 = "& Convert_SLV_To_Hex_String(conv5x_xi176_1159) & " elementx_x015x_xi174_1145 = "& Convert_SLV_To_Hex_String(elementx_x015x_xi174_1145) & " outputs:" & " addx_xi177_1164= "  & Convert_SLV_To_Hex_String(addx_xi177_1164));
      --
    end process; 
    -- binary operator OR_u64_u64_1163_inst
    process(conv5x_xi176_1159, elementx_x015x_xi174_1145) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi176_1159, elementx_x015x_xi174_1145, tmp_var);
      addx_xi177_1164 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u64_u64_613_inst flow-through 
    process(add_614) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:OR_u64_u64_613_inst:flowthrough inputs: " & " shl_602 = "& Convert_SLV_To_Hex_String(shl_602) & " conv24_609 = "& Convert_SLV_To_Hex_String(conv24_609) & " outputs:" & " add_614= "  & Convert_SLV_To_Hex_String(add_614));
      --
    end process; 
    -- binary operator OR_u64_u64_613_inst
    process(shl_602, conv24_609) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_602, conv24_609, tmp_var);
      add_614 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u64_u64_631_inst flow-through 
    process(add30_632) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:OR_u64_u64_631_inst:flowthrough inputs: " & " shl26_620 = "& Convert_SLV_To_Hex_String(shl26_620) & " conv29_627 = "& Convert_SLV_To_Hex_String(conv29_627) & " outputs:" & " add30_632= "  & Convert_SLV_To_Hex_String(add30_632));
      --
    end process; 
    -- binary operator OR_u64_u64_631_inst
    process(shl26_620, conv29_627) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl26_620, conv29_627, tmp_var);
      add30_632 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u64_u64_649_inst flow-through 
    process(add36_650) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:OR_u64_u64_649_inst:flowthrough inputs: " & " shl32_638 = "& Convert_SLV_To_Hex_String(shl32_638) & " conv35_645 = "& Convert_SLV_To_Hex_String(conv35_645) & " outputs:" & " add36_650= "  & Convert_SLV_To_Hex_String(add36_650));
      --
    end process; 
    -- binary operator OR_u64_u64_649_inst
    process(shl32_638, conv35_645) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl32_638, conv35_645, tmp_var);
      add36_650 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u64_u64_769_inst flow-through 
    process(addx_xi_770) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:OR_u64_u64_769_inst:flowthrough inputs: " & " conv5x_xi_765 = "& Convert_SLV_To_Hex_String(conv5x_xi_765) & " elementx_x015x_xi_751 = "& Convert_SLV_To_Hex_String(elementx_x015x_xi_751) & " outputs:" & " addx_xi_770= "  & Convert_SLV_To_Hex_String(addx_xi_770));
      --
    end process; 
    -- binary operator OR_u64_u64_769_inst
    process(conv5x_xi_765, elementx_x015x_xi_751) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi_765, elementx_x015x_xi_751, tmp_var);
      addx_xi_770 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_1008_inst flow-through 
    process(shl77_1009) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_1008_inst:flowthrough inputs: " & " add75_1003 = "& Convert_SLV_To_Hex_String(add75_1003) & " type_cast_1007_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1007_wire_constant) & " outputs:" & " shl77_1009= "  & Convert_SLV_To_Hex_String(shl77_1009));
      --
    end process; 
    -- binary operator SHL_u64_u64_1008_inst
    process(add75_1003) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add75_1003, type_cast_1007_wire_constant, tmp_var);
      shl77_1009 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_1026_inst flow-through 
    process(shl83_1027) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_1026_inst:flowthrough inputs: " & " add81_1021 = "& Convert_SLV_To_Hex_String(add81_1021) & " type_cast_1025_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1025_wire_constant) & " outputs:" & " shl83_1027= "  & Convert_SLV_To_Hex_String(shl83_1027));
      --
    end process; 
    -- binary operator SHL_u64_u64_1026_inst
    process(add81_1021) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add81_1021, type_cast_1025_wire_constant, tmp_var);
      shl83_1027 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_1073_inst flow-through 
    process(tmp237_1074) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_1073_inst:flowthrough inputs: " & " umax_1068 = "& Convert_SLV_To_Hex_String(umax_1068) & " type_cast_1072_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1072_wire_constant) & " outputs:" & " tmp237_1074= "  & Convert_SLV_To_Hex_String(tmp237_1074));
      --
    end process; 
    -- binary operator SHL_u64_u64_1073_inst
    process(umax_1068) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_1068, type_cast_1072_wire_constant, tmp_var);
      tmp237_1074 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_1169_inst flow-through 
    process(shlx_xi178_1170) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_1169_inst:flowthrough inputs: " & " addx_xi177_1164 = "& Convert_SLV_To_Hex_String(addx_xi177_1164) & " type_cast_1168_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1168_wire_constant) & " outputs:" & " shlx_xi178_1170= "  & Convert_SLV_To_Hex_String(shlx_xi178_1170));
      --
    end process; 
    -- binary operator SHL_u64_u64_1169_inst
    process(addx_xi177_1164) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi177_1164, type_cast_1168_wire_constant, tmp_var);
      shlx_xi178_1170 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_1198_inst flow-through 
    process(iNsTr_52_1199) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_1198_inst:flowthrough inputs: " & " mul58_862 = "& Convert_SLV_To_Hex_String(mul58_862) & " type_cast_1197_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1197_wire_constant) & " outputs:" & " iNsTr_52_1199= "  & Convert_SLV_To_Hex_String(iNsTr_52_1199));
      --
    end process; 
    -- binary operator SHL_u64_u64_1198_inst
    process(mul58_862) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul58_862, type_cast_1197_wire_constant, tmp_var);
      iNsTr_52_1199 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_1215_inst flow-through 
    process(shl12x_xi187_1216) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_1215_inst:flowthrough inputs: " & " shlx_xi178x_xlcssa_1189 = "& Convert_SLV_To_Hex_String(shlx_xi178x_xlcssa_1189) & " sh_promx_xi186_1211 = "& Convert_SLV_To_Hex_String(sh_promx_xi186_1211) & " outputs:" & " shl12x_xi187_1216= "  & Convert_SLV_To_Hex_String(shl12x_xi187_1216));
      --
    end process; 
    -- binary operator SHL_u64_u64_1215_inst
    process(shlx_xi178x_xlcssa_1189, sh_promx_xi186_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shlx_xi178x_xlcssa_1189, sh_promx_xi186_1211, tmp_var);
      shl12x_xi187_1216 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_486_inst flow-through 
    process(sext_487) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_486_inst:flowthrough inputs: " & " mul12_481 = "& Convert_SLV_To_Hex_String(mul12_481) & " type_cast_485_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_485_wire_constant) & " outputs:" & " sext_487= "  & Convert_SLV_To_Hex_String(sext_487));
      --
    end process; 
    -- binary operator SHL_u64_u64_486_inst
    process(mul12_481) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul12_481, type_cast_485_wire_constant, tmp_var);
      sext_487 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_601_inst flow-through 
    process(shl_602) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_601_inst:flowthrough inputs: " & " conv20_596 = "& Convert_SLV_To_Hex_String(conv20_596) & " type_cast_600_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_600_wire_constant) & " outputs:" & " shl_602= "  & Convert_SLV_To_Hex_String(shl_602));
      --
    end process; 
    -- binary operator SHL_u64_u64_601_inst
    process(conv20_596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv20_596, type_cast_600_wire_constant, tmp_var);
      shl_602 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_619_inst flow-through 
    process(shl26_620) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_619_inst:flowthrough inputs: " & " add_614 = "& Convert_SLV_To_Hex_String(add_614) & " type_cast_618_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_618_wire_constant) & " outputs:" & " shl26_620= "  & Convert_SLV_To_Hex_String(shl26_620));
      --
    end process; 
    -- binary operator SHL_u64_u64_619_inst
    process(add_614) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_614, type_cast_618_wire_constant, tmp_var);
      shl26_620 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_637_inst flow-through 
    process(shl32_638) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_637_inst:flowthrough inputs: " & " add30_632 = "& Convert_SLV_To_Hex_String(add30_632) & " type_cast_636_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_636_wire_constant) & " outputs:" & " shl32_638= "  & Convert_SLV_To_Hex_String(shl32_638));
      --
    end process; 
    -- binary operator SHL_u64_u64_637_inst
    process(add30_632) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add30_632, type_cast_636_wire_constant, tmp_var);
      shl32_638 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_684_inst flow-through 
    process(tmp253_685) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_684_inst:flowthrough inputs: " & " umax252_679 = "& Convert_SLV_To_Hex_String(umax252_679) & " type_cast_683_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_683_wire_constant) & " outputs:" & " tmp253_685= "  & Convert_SLV_To_Hex_String(tmp253_685));
      --
    end process; 
    -- binary operator SHL_u64_u64_684_inst
    process(umax252_679) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax252_679, type_cast_683_wire_constant, tmp_var);
      tmp253_685 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_775_inst flow-through 
    process(shlx_xi_776) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_775_inst:flowthrough inputs: " & " addx_xi_770 = "& Convert_SLV_To_Hex_String(addx_xi_770) & " type_cast_774_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_774_wire_constant) & " outputs:" & " shlx_xi_776= "  & Convert_SLV_To_Hex_String(shlx_xi_776));
      --
    end process; 
    -- binary operator SHL_u64_u64_775_inst
    process(addx_xi_770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_770, type_cast_774_wire_constant, tmp_var);
      shlx_xi_776 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_804_inst flow-through 
    process(iNsTr_38_805) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_804_inst:flowthrough inputs: " & " mul12_481 = "& Convert_SLV_To_Hex_String(mul12_481) & " type_cast_803_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_803_wire_constant) & " outputs:" & " iNsTr_38_805= "  & Convert_SLV_To_Hex_String(iNsTr_38_805));
      --
    end process; 
    -- binary operator SHL_u64_u64_804_inst
    process(mul12_481) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul12_481, type_cast_803_wire_constant, tmp_var);
      iNsTr_38_805 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_821_inst flow-through 
    process(shl12x_xi_822) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_821_inst:flowthrough inputs: " & " shlx_xix_xlcssa_795 = "& Convert_SLV_To_Hex_String(shlx_xix_xlcssa_795) & " sh_promx_xi_817 = "& Convert_SLV_To_Hex_String(sh_promx_xi_817) & " outputs:" & " shl12x_xi_822= "  & Convert_SLV_To_Hex_String(shl12x_xi_822));
      --
    end process; 
    -- binary operator SHL_u64_u64_821_inst
    process(shlx_xix_xlcssa_795, sh_promx_xi_817) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shlx_xix_xlcssa_795, sh_promx_xi_817, tmp_var);
      shl12x_xi_822 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_867_inst flow-through 
    process(sext171_868) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_867_inst:flowthrough inputs: " & " mul58_862 = "& Convert_SLV_To_Hex_String(mul58_862) & " type_cast_866_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_866_wire_constant) & " outputs:" & " sext171_868= "  & Convert_SLV_To_Hex_String(sext171_868));
      --
    end process; 
    -- binary operator SHL_u64_u64_867_inst
    process(mul58_862) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul58_862, type_cast_866_wire_constant, tmp_var);
      sext171_868 <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_990_inst flow-through 
    process(shl71_991) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SHL_u64_u64_990_inst:flowthrough inputs: " & " conv69_985 = "& Convert_SLV_To_Hex_String(conv69_985) & " type_cast_989_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_989_wire_constant) & " outputs:" & " shl71_991= "  & Convert_SLV_To_Hex_String(shl71_991));
      --
    end process; 
    -- binary operator SHL_u64_u64_990_inst
    process(conv69_985) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv69_985, type_cast_989_wire_constant, tmp_var);
      shl71_991 <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u64_u64_1369_inst flow-through 
    process(sub169_1370) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:SUB_u64_u64_1369_inst:flowthrough inputs: " & " conv165_1365 = "& Convert_SLV_To_Hex_String(conv165_1365) & " conv110_1357 = "& Convert_SLV_To_Hex_String(conv110_1357) & " outputs:" & " sub169_1370= "  & Convert_SLV_To_Hex_String(sub169_1370));
      --
    end process; 
    -- binary operator SUB_u64_u64_1369_inst
    process(conv165_1365, conv110_1357) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv165_1365, conv110_1357, tmp_var);
      sub169_1370 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u64_u1_502_inst flow-through 
    process(cmp195_503) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:UGT_u64_u1_502_inst:flowthrough inputs: " & " conv13_497 = "& Convert_SLV_To_Hex_String(conv13_497) & " type_cast_501_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_501_wire_constant) & " outputs:" & " cmp195_503= "  & Convert_SLV_To_Hex_String(cmp195_503));
      --
    end process; 
    -- binary operator UGT_u64_u1_502_inst
    process(conv13_497) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv13_497, type_cast_501_wire_constant, tmp_var);
      cmp195_503 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u64_u1_521_inst flow-through 
    process(tmp251_522) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:UGT_u64_u1_521_inst:flowthrough inputs: " & " tmp250_516 = "& Convert_SLV_To_Hex_String(tmp250_516) & " type_cast_520_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_520_wire_constant) & " outputs:" & " tmp251_522= "  & Convert_SLV_To_Hex_String(tmp251_522));
      --
    end process; 
    -- binary operator UGT_u64_u1_521_inst
    process(tmp250_516) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp250_516, type_cast_520_wire_constant, tmp_var);
      tmp251_522 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u64_u1_564_inst flow-through 
    process(tmp35_565) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:UGT_u64_u1_564_inst:flowthrough inputs: " & " tmp34_559 = "& Convert_SLV_To_Hex_String(tmp34_559) & " type_cast_563_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_563_wire_constant) & " outputs:" & " tmp35_565= "  & Convert_SLV_To_Hex_String(tmp35_565));
      --
    end process; 
    -- binary operator UGT_u64_u1_564_inst
    process(tmp34_559) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp34_559, type_cast_563_wire_constant, tmp_var);
      tmp35_565 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u64_u1_882_inst flow-through 
    process(cmp65191_883) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:UGT_u64_u1_882_inst:flowthrough inputs: " & " conv59_877 = "& Convert_SLV_To_Hex_String(conv59_877) & " type_cast_881_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_881_wire_constant) & " outputs:" & " cmp65191_883= "  & Convert_SLV_To_Hex_String(cmp65191_883));
      --
    end process; 
    -- binary operator UGT_u64_u1_882_inst
    process(conv59_877) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv59_877, type_cast_881_wire_constant, tmp_var);
      cmp65191_883 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u64_u1_901_inst flow-through 
    process(tmp236_902) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:UGT_u64_u1_901_inst:flowthrough inputs: " & " tmp235_896 = "& Convert_SLV_To_Hex_String(tmp235_896) & " type_cast_900_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_900_wire_constant) & " outputs:" & " tmp236_902= "  & Convert_SLV_To_Hex_String(tmp236_902));
      --
    end process; 
    -- binary operator UGT_u64_u1_901_inst
    process(tmp235_896) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp235_896, type_cast_900_wire_constant, tmp_var);
      tmp236_902 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u64_u1_953_inst flow-through 
    process(tmp24_954) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:UGT_u64_u1_953_inst:flowthrough inputs: " & " tmp23_948 = "& Convert_SLV_To_Hex_String(tmp23_948) & " type_cast_952_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_952_wire_constant) & " outputs:" & " tmp24_954= "  & Convert_SLV_To_Hex_String(tmp24_954));
      --
    end process; 
    -- binary operator UGT_u64_u1_953_inst
    process(tmp23_948) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp23_948, type_cast_952_wire_constant, tmp_var);
      tmp24_954 <= tmp_var; --
    end process;
    -- logger for split-operator XOR_u64_u64_1210_inst flow-through 
    process(sh_promx_xi186_1211) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:XOR_u64_u64_1210_inst:flowthrough inputs: " & " mulx_xi185_1205 = "& Convert_SLV_To_Hex_String(mulx_xi185_1205) & " type_cast_1209_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1209_wire_constant) & " outputs:" & " sh_promx_xi186_1211= "  & Convert_SLV_To_Hex_String(sh_promx_xi186_1211));
      --
    end process; 
    -- binary operator XOR_u64_u64_1210_inst
    process(mulx_xi185_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(mulx_xi185_1205, type_cast_1209_wire_constant, tmp_var);
      sh_promx_xi186_1211 <= tmp_var; --
    end process;
    -- logger for split-operator XOR_u64_u64_816_inst flow-through 
    process(sh_promx_xi_817) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:XOR_u64_u64_816_inst:flowthrough inputs: " & " mulx_xi_811 = "& Convert_SLV_To_Hex_String(mulx_xi_811) & " type_cast_815_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_815_wire_constant) & " outputs:" & " sh_promx_xi_817= "  & Convert_SLV_To_Hex_String(sh_promx_xi_817));
      --
    end process; 
    -- binary operator XOR_u64_u64_816_inst
    process(mulx_xi_811) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(mulx_xi_811, type_cast_815_wire_constant, tmp_var);
      sh_promx_xi_817 <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_1221_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1221_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_1221_index_offset:started:   inputs: " & " R_ix_x1x_xlcssa_1220_scaled = "& Convert_SLV_To_Hex_String(R_ix_x1x_xlcssa_1220_scaled) & " array_obj_ref_1221_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1221_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1221_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_1221_index_offset:finished:  outputs: " & " array_obj_ref_1221_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1221_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (82) : array_obj_ref_1221_index_offset 
    ApIntAdd_group_82: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_1220_scaled;
      array_obj_ref_1221_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1221_index_offset_req_0;
      array_obj_ref_1221_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1221_index_offset_req_1;
      array_obj_ref_1221_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_82_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_82_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_82",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 82
    -- logger for split-operator array_obj_ref_587_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_587_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_587_index_offset:started:   inputs: " & " R_indvar256_586_scaled = "& Convert_SLV_To_Hex_String(R_indvar256_586_scaled) & " array_obj_ref_587_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_587_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_587_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_587_index_offset:finished:  outputs: " & " array_obj_ref_587_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_587_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (83) : array_obj_ref_587_index_offset 
    ApIntAdd_group_83: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar256_586_scaled;
      array_obj_ref_587_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_587_index_offset_req_0;
      array_obj_ref_587_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_587_index_offset_req_1;
      array_obj_ref_587_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_83_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_83_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_83",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 83
    -- logger for split-operator array_obj_ref_827_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_827_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_827_index_offset:started:   inputs: " & " R_ix_x0x_xlcssa_826_scaled = "& Convert_SLV_To_Hex_String(R_ix_x0x_xlcssa_826_scaled) & " array_obj_ref_827_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_827_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_827_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_827_index_offset:finished:  outputs: " & " array_obj_ref_827_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_827_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (84) : array_obj_ref_827_index_offset 
    ApIntAdd_group_84: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_826_scaled;
      array_obj_ref_827_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_827_index_offset_req_0;
      array_obj_ref_827_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_827_index_offset_req_1;
      array_obj_ref_827_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_84_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_84_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_84",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 84
    -- logger for split-operator array_obj_ref_976_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_976_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_976_index_offset:started:   inputs: " & " R_indvar240_975_scaled = "& Convert_SLV_To_Hex_String(R_indvar240_975_scaled) & " array_obj_ref_976_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_976_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_976_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:array_obj_ref_976_index_offset:finished:  outputs: " & " array_obj_ref_976_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_976_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (85) : array_obj_ref_976_index_offset 
    ApIntAdd_group_85: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar240_975_scaled;
      array_obj_ref_976_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_976_index_offset_req_0;
      array_obj_ref_976_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_976_index_offset_req_1;
      array_obj_ref_976_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_85_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_85_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_85",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 85
    -- logger for split-operator type_cast_1355_inst flow-through 
    process(type_cast_1355_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1355_inst:flowthrough inputs: " & " call109_1232 = "& Convert_SLV_To_Hex_String(call109_1232) & " outputs:" & " type_cast_1355_wire= "  & Convert_SLV_To_Hex_String(type_cast_1355_wire));
      --
    end process; 
    -- unary operator type_cast_1355_inst
    process(call109_1232) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call109_1232, tmp_var);
      type_cast_1355_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1363_inst flow-through 
    process(type_cast_1363_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_1363_inst:flowthrough inputs: " & " call164_1360 = "& Convert_SLV_To_Hex_String(call164_1360) & " outputs:" & " type_cast_1363_wire= "  & Convert_SLV_To_Hex_String(type_cast_1363_wire));
      --
    end process; 
    -- unary operator type_cast_1363_inst
    process(call164_1360) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call164_1360, tmp_var);
      type_cast_1363_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_551_inst flow-through 
    process(type_cast_551_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_551_inst:flowthrough inputs: " & " tmp32_548 = "& Convert_SLV_To_Hex_String(tmp32_548) & " outputs:" & " type_cast_551_wire= "  & Convert_SLV_To_Hex_String(type_cast_551_wire));
      --
    end process; 
    -- unary operator type_cast_551_inst
    process(tmp32_548) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp32_548, tmp_var);
      type_cast_551_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_940_inst flow-through 
    process(type_cast_940_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:type_cast_940_inst:flowthrough inputs: " & " tmp21_937 = "& Convert_SLV_To_Hex_String(tmp21_937) & " outputs:" & " type_cast_940_wire= "  & Convert_SLV_To_Hex_String(type_cast_940_wire));
      --
    end process; 
    -- unary operator type_cast_940_inst
    process(tmp21_937) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp21_937, tmp_var);
      type_cast_940_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator ptr_deref_1225_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1225_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_1225_store_0:started:   inputs: " & " ptr_deref_1225_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1225_word_address_0) & " ptr_deref_1225_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1225_data_0));
          --
        end if; 
        if ptr_deref_1225_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_1225_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_1041_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1041_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_1041_store_0:started:   inputs: " & " ptr_deref_1041_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1041_word_address_0) & " ptr_deref_1041_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1041_data_0));
          --
        end if; 
        if ptr_deref_1041_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_1041_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1225_store_0_req_0,
      ptr_deref_1225_store_0_ack_0,
      ptr_deref_1225_store_0_req_1,
      ptr_deref_1225_store_0_ack_1,
      "ptr_deref_1225_store_0",
      "memory_space_0" ,
      ptr_deref_1225_data_0,
      ptr_deref_1225_word_address_0,
      "ptr_deref_1225_data_0",
      "ptr_deref_1225_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1041_store_0_req_0,
      ptr_deref_1041_store_0_ack_0,
      ptr_deref_1041_store_0_req_1,
      ptr_deref_1041_store_0_ack_1,
      "ptr_deref_1041_store_0",
      "memory_space_0" ,
      ptr_deref_1041_data_0,
      ptr_deref_1041_word_address_0,
      "ptr_deref_1041_data_0",
      "ptr_deref_1041_word_address_0" -- 
    );
    -- shared store operator group (0) : ptr_deref_1225_store_0 ptr_deref_1041_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1225_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1041_store_0_req_0;
      ptr_deref_1225_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1041_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1225_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1041_store_0_req_1;
      ptr_deref_1225_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1041_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1225_word_address_0 & ptr_deref_1041_word_address_0;
      data_in <= ptr_deref_1225_data_0 & ptr_deref_1041_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logger for split-operator ptr_deref_652_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_652_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_652_store_0:started:   inputs: " & " ptr_deref_652_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_652_word_address_0) & " ptr_deref_652_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_652_data_0));
          --
        end if; 
        if ptr_deref_652_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_652_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_831_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_831_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_831_store_0:started:   inputs: " & " ptr_deref_831_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_831_word_address_0) & " ptr_deref_831_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_831_data_0));
          --
        end if; 
        if ptr_deref_831_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:ptr_deref_831_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_652_store_0_req_0,
      ptr_deref_652_store_0_ack_0,
      ptr_deref_652_store_0_req_1,
      ptr_deref_652_store_0_ack_1,
      "ptr_deref_652_store_0",
      "memory_space_1" ,
      ptr_deref_652_data_0,
      ptr_deref_652_word_address_0,
      "ptr_deref_652_data_0",
      "ptr_deref_652_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_831_store_0_req_0,
      ptr_deref_831_store_0_ack_0,
      ptr_deref_831_store_0_req_1,
      ptr_deref_831_store_0_ack_1,
      "ptr_deref_831_store_0",
      "memory_space_1" ,
      ptr_deref_831_data_0,
      ptr_deref_831_word_address_0,
      "ptr_deref_831_data_0",
      "ptr_deref_831_word_address_0" -- 
    );
    -- shared store operator group (1) : ptr_deref_652_store_0 ptr_deref_831_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_652_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_831_store_0_req_0;
      ptr_deref_652_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_831_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_652_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_831_store_0_req_1;
      ptr_deref_652_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_831_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_652_word_address_0 & ptr_deref_831_word_address_0;
      data_in <= ptr_deref_652_data_0 & ptr_deref_831_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- logger for split-operator RPIPE_maxpool_input_pipe_443_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_443_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_443_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_443_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_443_inst:finished:  outputs: " & " call2_444= "  & Convert_SLV_To_Hex_String(call2_444));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_455_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_455_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_455_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_455_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_455_inst:finished:  outputs: " & " call6_456= "  & Convert_SLV_To_Hex_String(call6_456));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_458_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_458_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_458_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_458_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_458_inst:finished:  outputs: " & " call7_459= "  & Convert_SLV_To_Hex_String(call7_459));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_760_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_760_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_760_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_760_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_760_inst:finished:  outputs: " & " callx_xi_761= "  & Convert_SLV_To_Hex_String(callx_xi_761));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_640_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_640_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_640_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_640_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_640_inst:finished:  outputs: " & " call33_641= "  & Convert_SLV_To_Hex_String(call33_641));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_622_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_622_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_622_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_622_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_622_inst:finished:  outputs: " & " call27_623= "  & Convert_SLV_To_Hex_String(call27_623));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_446_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_446_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_446_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_446_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_446_inst:finished:  outputs: " & " call3_447= "  & Convert_SLV_To_Hex_String(call3_447));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_591_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_591_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_591_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_591_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_591_inst:finished:  outputs: " & " call19_592= "  & Convert_SLV_To_Hex_String(call19_592));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_604_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_604_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_604_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_604_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_604_inst:finished:  outputs: " & " call22_605= "  & Convert_SLV_To_Hex_String(call22_605));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_440_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_440_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_440_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_440_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_440_inst:finished:  outputs: " & " call1_441= "  & Convert_SLV_To_Hex_String(call1_441));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_452_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_452_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_452_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_452_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_452_inst:finished:  outputs: " & " call5_453= "  & Convert_SLV_To_Hex_String(call5_453));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_449_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_449_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_449_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_449_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_449_inst:finished:  outputs: " & " call4_450= "  & Convert_SLV_To_Hex_String(call4_450));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_437_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_437_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_437_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_437_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_437_inst:finished:  outputs: " & " call_438= "  & Convert_SLV_To_Hex_String(call_438));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_980_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_980_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_980_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_980_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_980_inst:finished:  outputs: " & " call68_981= "  & Convert_SLV_To_Hex_String(call68_981));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_993_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_993_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_993_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_993_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_993_inst:finished:  outputs: " & " call72_994= "  & Convert_SLV_To_Hex_String(call72_994));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_1011_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_1011_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_1011_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_1011_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_1011_inst:finished:  outputs: " & " call78_1012= "  & Convert_SLV_To_Hex_String(call78_1012));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_1029_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_1029_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_1029_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_1029_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_1029_inst:finished:  outputs: " & " call84_1030= "  & Convert_SLV_To_Hex_String(call84_1030));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_1154_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_1154_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_1154_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_1154_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:RPIPE_maxpool_input_pipe_1154_inst:finished:  outputs: " & " callx_xi175_1155= "  & Convert_SLV_To_Hex_String(callx_xi175_1155));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_443_inst RPIPE_maxpool_input_pipe_455_inst RPIPE_maxpool_input_pipe_458_inst RPIPE_maxpool_input_pipe_760_inst RPIPE_maxpool_input_pipe_640_inst RPIPE_maxpool_input_pipe_622_inst RPIPE_maxpool_input_pipe_446_inst RPIPE_maxpool_input_pipe_591_inst RPIPE_maxpool_input_pipe_604_inst RPIPE_maxpool_input_pipe_440_inst RPIPE_maxpool_input_pipe_452_inst RPIPE_maxpool_input_pipe_449_inst RPIPE_maxpool_input_pipe_437_inst RPIPE_maxpool_input_pipe_980_inst RPIPE_maxpool_input_pipe_993_inst RPIPE_maxpool_input_pipe_1011_inst RPIPE_maxpool_input_pipe_1029_inst RPIPE_maxpool_input_pipe_1154_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(287 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 17 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 17 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 17 downto 0);
      signal guard_vector : std_logic_vector( 17 downto 0);
      constant outBUFs : IntegerArray(17 downto 0) := (17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(17 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false);
      constant guardBuffering: IntegerArray(17 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2);
      -- 
    begin -- 
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_443_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_455_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_458_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_760_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_640_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_622_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_446_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_591_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_604_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_440_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_452_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_449_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_437_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_980_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_993_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_1011_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_1029_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1154_inst_req_0;
      RPIPE_maxpool_input_pipe_443_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_455_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_458_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_760_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_640_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_622_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_446_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_591_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_604_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_440_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_452_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_449_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_437_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_980_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_993_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_1011_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_1029_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1154_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_443_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_455_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_458_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_760_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_640_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_622_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_446_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_591_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_604_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_440_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_452_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_449_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_437_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_980_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_993_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_1011_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_1029_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1154_inst_req_1;
      RPIPE_maxpool_input_pipe_443_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_455_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_458_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_760_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_640_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_622_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_446_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_591_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_604_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_440_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_452_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_449_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_437_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_980_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_993_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_1011_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_1029_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1154_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      call2_444 <= data_out(287 downto 272);
      call6_456 <= data_out(271 downto 256);
      call7_459 <= data_out(255 downto 240);
      callx_xi_761 <= data_out(239 downto 224);
      call33_641 <= data_out(223 downto 208);
      call27_623 <= data_out(207 downto 192);
      call3_447 <= data_out(191 downto 176);
      call19_592 <= data_out(175 downto 160);
      call22_605 <= data_out(159 downto 144);
      call1_441 <= data_out(143 downto 128);
      call5_453 <= data_out(127 downto 112);
      call4_450 <= data_out(111 downto 96);
      call_438 <= data_out(95 downto 80);
      call68_981 <= data_out(79 downto 64);
      call72_994 <= data_out(63 downto 48);
      call78_1012 <= data_out(47 downto 32);
      call84_1030 <= data_out(31 downto 16);
      callx_xi175_1155 <= data_out(15 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 18, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 16,  num_reqs => 18,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_elapsed_time_pipe_1371_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_elapsed_time_pipe_1371_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:WPIPE_elapsed_time_pipe_1371_inst:started:   PipeWrite to elapsed_time_pipe inputs: " & " sub169_1370 = "& Convert_SLV_To_Hex_String(sub169_1370));
          --
        end if; 
        if WPIPE_elapsed_time_pipe_1371_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:WPIPE_elapsed_time_pipe_1371_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_elapsed_time_pipe_1371_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1371_inst_req_0;
      WPIPE_elapsed_time_pipe_1371_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1371_inst_req_1;
      WPIPE_elapsed_time_pipe_1371_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub169_1370;
      elapsed_time_pipe_write_0_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator WPIPE_maxpool_output_pipe_1247_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_maxpool_output_pipe_1247_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:WPIPE_maxpool_output_pipe_1247_inst:started:   PipeWrite to maxpool_output_pipe inputs: " & " type_cast_1249_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1249_wire_constant));
          --
        end if; 
        if WPIPE_maxpool_output_pipe_1247_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:WPIPE_maxpool_output_pipe_1247_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (1) : WPIPE_maxpool_output_pipe_1247_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1247_inst_req_0;
      WPIPE_maxpool_output_pipe_1247_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1247_inst_req_1;
      WPIPE_maxpool_output_pipe_1247_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1249_wire_constant;
      maxpool_output_pipe_write_1_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logger for split-operator WPIPE_num_out_pipe_1244_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_num_out_pipe_1244_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:WPIPE_num_out_pipe_1244_inst:started:   PipeWrite to num_out_pipe inputs: " & " mul129_1243 = "& Convert_SLV_To_Hex_String(mul129_1243));
          --
        end if; 
        if WPIPE_num_out_pipe_1244_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:WPIPE_num_out_pipe_1244_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (2) : WPIPE_num_out_pipe_1244_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_1244_inst_req_0;
      WPIPE_num_out_pipe_1244_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_num_out_pipe_1244_inst_req_1;
      WPIPE_num_out_pipe_1244_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= mul129_1243;
      num_out_pipe_write_2_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- logger for split-operator call_stmt_1360_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1360_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:call_stmt_1360_call:started:  Call to module timer inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if call_stmt_1360_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:call_stmt_1360_call:finished:  outputs: " & " call164_1360= "  & Convert_SLV_To_Hex_String(call164_1360));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_1232_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1232_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:call_stmt_1232_call:started:  Call to module timer inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if call_stmt_1232_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:call_stmt_1232_call:finished:  outputs: " & " call109_1232= "  & Convert_SLV_To_Hex_String(call109_1232));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_1360_call call_stmt_1232_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1360_call_req_0;
      reqL_unguarded(0) <= call_stmt_1232_call_req_0;
      call_stmt_1360_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1232_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1360_call_req_1;
      reqR_unguarded(0) <= call_stmt_1232_call_req_1;
      call_stmt_1360_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1232_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call164_1360 <= data_out(127 downto 64);
      call109_1232 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_1327_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1327_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:call_stmt_1327_call:started:  Call to module loadKernelChannel inputs: " & " conv135_1320 = "& Convert_SLV_To_Hex_String(conv135_1320) & " conv141_1324 = "& Convert_SLV_To_Hex_String(conv141_1324));
          --
        end if; 
        if call_stmt_1327_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:call_stmt_1327_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_1327_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1327_call_req_0;
      call_stmt_1327_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1327_call_req_1;
      call_stmt_1327_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv135_1320 & conv141_1324;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 128,
        owidth => 128,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(127 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- logger for split-operator call_stmt_1334_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1334_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:call_stmt_1334_call:started:  Call to module access_T inputs: " & " mul116_1238 = "& Convert_SLV_To_Hex_String(mul116_1238) & " call3_447 = "& Convert_SLV_To_Hex_String(call3_447) & " sub_1256 = "& Convert_SLV_To_Hex_String(sub_1256) & " sub149_1262 = "& Convert_SLV_To_Hex_String(sub149_1262) & " call2_444 = "& Convert_SLV_To_Hex_String(call2_444) & " call1_441 = "& Convert_SLV_To_Hex_String(call1_441));
          --
        end if; 
        if call_stmt_1334_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolution3D:DP:call_stmt_1334_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (2) : call_stmt_1334_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1334_call_req_0;
      call_stmt_1334_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1334_call_req_1;
      call_stmt_1334_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul116_1238 & call3_447 & sub_1256 & sub149_1262 & call2_444 & call1_441;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 96,
        owidth => 96,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(95 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_3268_start: Boolean;
  signal convolve_CP_3268_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_kernel_pipe1_1469_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1494_inst_ack_0 : boolean;
  signal nacc_1454_1405_buf_req_0 : boolean;
  signal n_out_count_1483_1410_buf_ack_0 : boolean;
  signal WPIPE_input_done_pipe_1490_inst_req_0 : boolean;
  signal SUB_u32_u32_1435_inst_req_1 : boolean;
  signal n_out_count_1483_1410_buf_req_0 : boolean;
  signal type_cast_1496_inst_ack_1 : boolean;
  signal type_cast_1496_inst_req_1 : boolean;
  signal RPIPE_input_pipe1_1413_inst_ack_1 : boolean;
  signal WPIPE_input_done_pipe_1490_inst_ack_1 : boolean;
  signal RPIPE_input_pipe1_1413_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1494_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_1490_inst_req_1 : boolean;
  signal type_cast_1496_inst_ack_0 : boolean;
  signal n_out_count_1483_1410_buf_ack_1 : boolean;
  signal RPIPE_input_pipe1_1413_inst_ack_0 : boolean;
  signal RPIPE_input_pipe1_1413_inst_req_0 : boolean;
  signal nacc_1454_1405_buf_ack_0 : boolean;
  signal phi_stmt_1406_ack_0 : boolean;
  signal SUB_u32_u32_1435_inst_ack_0 : boolean;
  signal SUB_u32_u32_1435_inst_req_0 : boolean;
  signal nacc_1454_1405_buf_ack_1 : boolean;
  signal nacc_1454_1405_buf_req_1 : boolean;
  signal WPIPE_kernel_pipe1_1469_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_1469_inst_req_1 : boolean;
  signal n_out_count_1483_1410_buf_req_1 : boolean;
  signal phi_stmt_1406_req_0 : boolean;
  signal RPIPE_kernel_pipe1_1421_inst_ack_1 : boolean;
  signal WPIPE_input_done_pipe_1490_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_1421_inst_req_1 : boolean;
  signal type_cast_1496_inst_req_0 : boolean;
  signal phi_stmt_1406_req_1 : boolean;
  signal do_while_stmt_1396_branch_ack_1 : boolean;
  signal SUB_u32_u32_1435_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe1_1421_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe1_1469_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_1421_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1494_inst_req_1 : boolean;
  signal do_while_stmt_1396_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1494_inst_ack_1 : boolean;
  signal RPIPE_num_out_pipe_1382_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1382_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1382_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_1382_inst_ack_1 : boolean;
  signal RPIPE_size_pipe_1385_inst_req_0 : boolean;
  signal RPIPE_size_pipe_1385_inst_ack_0 : boolean;
  signal RPIPE_size_pipe_1385_inst_req_1 : boolean;
  signal RPIPE_size_pipe_1385_inst_ack_1 : boolean;
  signal do_while_stmt_1396_branch_req_0 : boolean;
  signal phi_stmt_1398_req_1 : boolean;
  signal phi_stmt_1398_req_0 : boolean;
  signal phi_stmt_1398_ack_0 : boolean;
  signal nmycount_1462_1401_buf_req_0 : boolean;
  signal nmycount_1462_1401_buf_ack_0 : boolean;
  signal nmycount_1462_1401_buf_req_1 : boolean;
  signal nmycount_1462_1401_buf_ack_1 : boolean;
  signal phi_stmt_1402_req_1 : boolean;
  signal phi_stmt_1402_req_0 : boolean;
  signal phi_stmt_1402_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_3268_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_3268_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_3268_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_3268_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,convolve_CP_3268_start,"convolve cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,convolve_CP_3268_symbol, "convolve cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_3268: Block -- control-path 
    signal convolve_CP_3268_elements: BooleanArray(104 downto 0);
    -- 
  begin -- 
    convolve_CP_3268_elements(0) <= convolve_CP_3268_start;
    convolve_CP_3268_symbol <= convolve_CP_3268_elements(1);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1380/$entry
      -- CP-element group 0: 	 branch_block_stmt_1380/branch_block_stmt_1380__entry__
      -- CP-element group 0: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395__entry__
      -- CP-element group 0: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/$entry
      -- CP-element group 0: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_num_out_pipe_1382_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_num_out_pipe_1382_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_num_out_pipe_1382_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_size_pipe_1385_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_size_pipe_1385_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_size_pipe_1385_Sample/rr
      -- 
    -- logger for CP element group convolve_CP_3268_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_num_out_pipe_1382_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_size_pipe_1385_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(0), ack => RPIPE_num_out_pipe_1382_inst_req_0); -- 
    rr_3304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(0), ack => RPIPE_size_pipe_1385_inst_req_0); -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	104 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1380/$exit
      -- CP-element group 1: 	 branch_block_stmt_1380/branch_block_stmt_1380__exit__
      -- CP-element group 1: 	 branch_block_stmt_1380/do_while_stmt_1396__exit__
      -- 
    -- logger for CP element group convolve_CP_3268_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(1) <= convolve_CP_3268_elements(104);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_num_out_pipe_1382_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_num_out_pipe_1382_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_num_out_pipe_1382_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_num_out_pipe_1382_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_num_out_pipe_1382_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_num_out_pipe_1382_Update/cr
      -- 
    -- logger for CP element group convolve_CP_3268_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_num_out_pipe_1382_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_num_out_pipe_1382_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_3291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1382_inst_ack_0, ack => convolve_CP_3268_elements(2)); -- 
    cr_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(2), ack => RPIPE_num_out_pipe_1382_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_num_out_pipe_1382_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_num_out_pipe_1382_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_num_out_pipe_1382_Update/ca
      -- 
    -- logger for CP element group convolve_CP_3268_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_num_out_pipe_1382_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1382_inst_ack_1, ack => convolve_CP_3268_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_size_pipe_1385_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_size_pipe_1385_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_size_pipe_1385_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_size_pipe_1385_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_size_pipe_1385_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_size_pipe_1385_Update/cr
      -- 
    -- logger for CP element group convolve_CP_3268_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_size_pipe_1385_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_size_pipe_1385_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_3305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1385_inst_ack_0, ack => convolve_CP_3268_elements(4)); -- 
    cr_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(4), ack => RPIPE_size_pipe_1385_inst_req_1); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_size_pipe_1385_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_size_pipe_1385_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/RPIPE_size_pipe_1385_Update/ca
      -- 
    -- logger for CP element group convolve_CP_3268_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_size_pipe_1385_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1385_inst_ack_1, ack => convolve_CP_3268_elements(5)); -- 
    -- CP-element group 6:  join  transition  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395__exit__
      -- CP-element group 6: 	 branch_block_stmt_1380/do_while_stmt_1396__entry__
      -- CP-element group 6: 	 branch_block_stmt_1380/assign_stmt_1383_to_assign_stmt_1395/$exit
      -- 
    -- logger for CP element group convolve_CP_3268_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    convolve_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "convolve_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(3) & convolve_CP_3268_elements(5);
      gj_convolve_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1380/do_while_stmt_1396/$entry
      -- CP-element group 7: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396__entry__
      -- 
    -- logger for CP element group convolve_CP_3268_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(7) <= convolve_CP_3268_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	104 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396__exit__
      -- 
    -- logger for CP element group convolve_CP_3268_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1380/do_while_stmt_1396/loop_back
      -- 
    -- logger for CP element group convolve_CP_3268_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	102 
    -- CP-element group 10: 	103 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1380/do_while_stmt_1396/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_1380/do_while_stmt_1396/loop_taken/$entry
      -- CP-element group 10: 	 branch_block_stmt_1380/do_while_stmt_1396/condition_done
      -- 
    -- logger for CP element group convolve_CP_3268_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(10) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(10) <= convolve_CP_3268_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	101 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1380/do_while_stmt_1396/loop_body_done
      -- 
    -- logger for CP element group convolve_CP_3268_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(11) <= convolve_CP_3268_elements(101);
    -- CP-element group 12:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	24 
    -- CP-element group 12: 	43 
    -- CP-element group 12: 	62 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group convolve_CP_3268_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(12) <= convolve_CP_3268_elements(9);
    -- CP-element group 13:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	26 
    -- CP-element group 13: 	45 
    -- CP-element group 13: 	64 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group convolve_CP_3268_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(13) <= convolve_CP_3268_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	21 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	38 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	57 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	79 
    -- CP-element group 14: 	83 
    -- CP-element group 14: 	100 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/loop_body_start
      -- 
    -- logger for CP element group convolve_CP_3268_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	100 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/condition_evaluated
      -- 
    -- logger for CP element group convolve_CP_3268_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:do_while_stmt_1396_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_3325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(15), ack => do_while_stmt_1396_branch_req_0); -- 
    convolve_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(19) & convolve_CP_3268_elements(100);
      gj_convolve_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	37 
    -- CP-element group 16: 	56 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	39 
    -- CP-element group 16: 	58 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/aggregated_phi_sample_req
      -- CP-element group 16: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_sample_start__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    convolve_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(20) & convolve_CP_3268_elements(37) & convolve_CP_3268_elements(56) & convolve_CP_3268_elements(19);
      gj_convolve_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	22 
    -- CP-element group 17: 	40 
    -- CP-element group 17: 	59 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	76 
    -- CP-element group 17: 	80 
    -- CP-element group 17: 	84 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	37 
    -- CP-element group 17: 	56 
    -- CP-element group 17:  members (4) 
      -- CP-element group 17: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/aggregated_phi_sample_ack
      -- CP-element group 17: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_sample_completed_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    convolve_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(22) & convolve_CP_3268_elements(40) & convolve_CP_3268_elements(59);
      gj_convolve_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: 	38 
    -- CP-element group 18: 	57 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	60 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/aggregated_phi_update_req
      -- CP-element group 18: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_update_start__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    convolve_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(21) & convolve_CP_3268_elements(38) & convolve_CP_3268_elements(57);
      gj_convolve_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	42 
    -- CP-element group 19: 	61 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group convolve_CP_3268_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    convolve_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(23) & convolve_CP_3268_elements(42) & convolve_CP_3268_elements(61);
      gj_convolve_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: 	86 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_sample_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(20) fired."); 
        -- 
      end if; --
    end process; 
    convolve_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(14) & convolve_CP_3268_elements(17) & convolve_CP_3268_elements(86);
      gj_convolve_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	14 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	91 
    -- CP-element group 21: 	95 
    -- CP-element group 21: 	98 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_update_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    convolve_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(14) & convolve_CP_3268_elements(91) & convolve_CP_3268_elements(95) & convolve_CP_3268_elements(98);
      gj_convolve_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	17 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_sample_completed__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(22) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: 	90 
    -- CP-element group 23: 	93 
    -- CP-element group 23: 	97 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_update_completed__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(23) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	12 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_loopback_trigger
      -- 
    -- logger for CP element group convolve_CP_3268_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(24) <= convolve_CP_3268_elements(12);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_loopback_sample_req
      -- CP-element group 25: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_loopback_sample_req_ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:phi_stmt_1398_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1398_loopback_sample_req_3340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1398_loopback_sample_req_3340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(25), ack => phi_stmt_1398_req_1); -- 
    -- Element group convolve_CP_3268_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	13 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_entry_trigger
      -- 
    -- logger for CP element group convolve_CP_3268_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(26) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(26) <= convolve_CP_3268_elements(13);
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_entry_sample_req
      -- CP-element group 27: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_entry_sample_req_ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:phi_stmt_1398_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1398_entry_sample_req_3343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1398_entry_sample_req_3343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(27), ack => phi_stmt_1398_req_0); -- 
    -- Element group convolve_CP_3268_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_phi_mux_ack
      -- CP-element group 28: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1398_phi_mux_ack_ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:phi_stmt_1398_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1398_phi_mux_ack_3346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1398_ack_0, ack => convolve_CP_3268_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_mcount_var_1400_sample_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_mcount_var_1400_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_mcount_var_1400_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_mcount_var_1400_sample_completed_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(29) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_mcount_var_1400_update_start__ps
      -- CP-element group 30: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_mcount_var_1400_update_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(30) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_mcount_var_1400_update_completed__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(31) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(31) <= convolve_CP_3268_elements(32);
    -- CP-element group 32:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	31 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_mcount_var_1400_update_completed_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(32) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(32) is a control-delay.
    cp_element_32_delay: control_delay_element  generic map(name => " 32_delay", delay_value => 1)  port map(req => convolve_CP_3268_elements(30), ack => convolve_CP_3268_elements(32), clk => clk, reset =>reset);
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_Sample/req
      -- 
    -- logger for CP element group convolve_CP_3268_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:nmycount_1462_1401_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(33), ack => nmycount_1462_1401_buf_req_0); -- 
    -- Element group convolve_CP_3268_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_update_start__ps
      -- CP-element group 34: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_Update/req
      -- 
    -- logger for CP element group convolve_CP_3268_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:nmycount_1462_1401_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(34), ack => nmycount_1462_1401_buf_req_1); -- 
    -- Element group convolve_CP_3268_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_Sample/ack
      -- 
    -- logger for CP element group convolve_CP_3268_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:nmycount_1462_1401_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1462_1401_buf_ack_0, ack => convolve_CP_3268_elements(35)); -- 
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nmycount_1401_Update/ack
      -- 
    -- logger for CP element group convolve_CP_3268_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:nmycount_1462_1401_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1462_1401_buf_ack_1, ack => convolve_CP_3268_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	17 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	82 
    -- CP-element group 37: 	86 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	16 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_sample_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(37) fired."); 
        -- 
      end if; --
    end process; 
    convolve_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(14) & convolve_CP_3268_elements(17) & convolve_CP_3268_elements(78) & convolve_CP_3268_elements(82) & convolve_CP_3268_elements(86);
      gj_convolve_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	14 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	95 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	18 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_update_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(38) fired."); 
        -- 
      end if; --
    end process; 
    convolve_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(14) & convolve_CP_3268_elements(95);
      gj_convolve_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	16 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_sample_start__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(39) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(39) <= convolve_CP_3268_elements(16);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	17 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_sample_completed__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(40) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_update_start__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(41) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(41) <= convolve_CP_3268_elements(18);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	19 
    -- CP-element group 42: 	93 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_update_completed__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(42) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	12 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_loopback_trigger
      -- 
    -- logger for CP element group convolve_CP_3268_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(43) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(43) <= convolve_CP_3268_elements(12);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_loopback_sample_req_ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:phi_stmt_1402_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1402_loopback_sample_req_3384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1402_loopback_sample_req_3384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(44), ack => phi_stmt_1402_req_1); -- 
    -- Element group convolve_CP_3268_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	13 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_entry_trigger
      -- 
    -- logger for CP element group convolve_CP_3268_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(45) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(45) <= convolve_CP_3268_elements(13);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_entry_sample_req_ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:phi_stmt_1402_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1402_entry_sample_req_3387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1402_entry_sample_req_3387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(46), ack => phi_stmt_1402_req_0); -- 
    -- Element group convolve_CP_3268_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1402_phi_mux_ack_ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:phi_stmt_1402_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1402_phi_mux_ack_3390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1402_ack_0, ack => convolve_CP_3268_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_acc_var_1404_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_acc_var_1404_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_acc_var_1404_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_acc_var_1404_sample_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(48) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_acc_var_1404_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_acc_var_1404_update_start__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(49) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_acc_var_1404_update_completed__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(50) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(50) <= convolve_CP_3268_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_acc_var_1404_update_completed_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(51) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => convolve_CP_3268_elements(49), ack => convolve_CP_3268_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_Sample/$entry
      -- 
    -- logger for CP element group convolve_CP_3268_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:nacc_1454_1405_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(52), ack => nacc_1454_1405_buf_req_0); -- 
    -- Element group convolve_CP_3268_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_Update/req
      -- CP-element group 53: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_update_start_
      -- CP-element group 53: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_update_start__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:nacc_1454_1405_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(53), ack => nacc_1454_1405_buf_req_1); -- 
    -- Element group convolve_CP_3268_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_Sample/$exit
      -- 
    -- logger for CP element group convolve_CP_3268_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:nacc_1454_1405_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1454_1405_buf_ack_0, ack => convolve_CP_3268_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_nacc_1405_update_completed_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:nacc_1454_1405_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1454_1405_buf_ack_1, ack => convolve_CP_3268_elements(55)); -- 
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	14 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	17 
    -- CP-element group 56: 	86 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	16 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_sample_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(56) fired."); 
        -- 
      end if; --
    end process; 
    convolve_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(14) & convolve_CP_3268_elements(17) & convolve_CP_3268_elements(86);
      gj_convolve_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	14 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	88 
    -- CP-element group 57: 	91 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	18 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_update_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(57) fired."); 
        -- 
      end if; --
    end process; 
    convolve_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(14) & convolve_CP_3268_elements(88) & convolve_CP_3268_elements(91);
      gj_convolve_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	16 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_sample_start__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(58) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(58) <= convolve_CP_3268_elements(16);
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	17 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_sample_completed__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(59) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	18 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_update_start__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(60) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(60) <= convolve_CP_3268_elements(18);
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	19 
    -- CP-element group 61: 	87 
    -- CP-element group 61: 	90 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_update_completed__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(61) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(61) is bound as output of CP function.
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	12 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_loopback_trigger
      -- 
    -- logger for CP element group convolve_CP_3268_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(62) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(62) <= convolve_CP_3268_elements(12);
    -- CP-element group 63:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_loopback_sample_req_ps
      -- CP-element group 63: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_loopback_sample_req
      -- 
    -- logger for CP element group convolve_CP_3268_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:phi_stmt_1406_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1406_loopback_sample_req_3428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1406_loopback_sample_req_3428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(63), ack => phi_stmt_1406_req_1); -- 
    -- Element group convolve_CP_3268_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	13 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_entry_trigger
      -- 
    -- logger for CP element group convolve_CP_3268_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(64) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(64) <= convolve_CP_3268_elements(13);
    -- CP-element group 65:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_entry_sample_req
      -- CP-element group 65: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_entry_sample_req_ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:phi_stmt_1406_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1406_entry_sample_req_3431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1406_entry_sample_req_3431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(65), ack => phi_stmt_1406_req_0); -- 
    -- Element group convolve_CP_3268_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_phi_mux_ack_ps
      -- CP-element group 66: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/phi_stmt_1406_phi_mux_ack
      -- 
    -- logger for CP element group convolve_CP_3268_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:phi_stmt_1406_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1406_phi_mux_ack_3434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1406_ack_0, ack => convolve_CP_3268_elements(66)); -- 
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1409_sample_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1409_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1409_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1409_sample_completed__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(67) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1409_update_start_
      -- CP-element group 68: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1409_update_start__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(68) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1409_update_completed__ps
      -- 
    -- logger for CP element group convolve_CP_3268_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(69) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(69) <= convolve_CP_3268_elements(70);
    -- CP-element group 70:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	69 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1409_update_completed_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(70) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => convolve_CP_3268_elements(68), ack => convolve_CP_3268_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_sample_start__ps
      -- CP-element group 71: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_sample_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(71) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:n_out_count_1483_1410_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(71), ack => n_out_count_1483_1410_buf_req_0); -- 
    -- Element group convolve_CP_3268_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_update_start__ps
      -- CP-element group 72: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_Update/req
      -- CP-element group 72: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_update_start_
      -- CP-element group 72: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_Update/$entry
      -- 
    -- logger for CP element group convolve_CP_3268_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(72) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:n_out_count_1483_1410_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(72), ack => n_out_count_1483_1410_buf_req_1); -- 
    -- Element group convolve_CP_3268_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_sample_completed__ps
      -- CP-element group 73: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_sample_completed_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:n_out_count_1483_1410_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1483_1410_buf_ack_0, ack => convolve_CP_3268_elements(73)); -- 
    -- CP-element group 74:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_update_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/R_n_out_count_1410_update_completed_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:n_out_count_1483_1410_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1483_1410_buf_ack_1, ack => convolve_CP_3268_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	78 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_input_pipe1_1413_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_input_pipe1_1413_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_input_pipe1_1413_sample_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_input_pipe1_1413_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(75), ack => RPIPE_input_pipe1_1413_inst_req_0); -- 
    convolve_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(14) & convolve_CP_3268_elements(78);
      gj_convolve_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	17 
    -- CP-element group 76: 	77 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	95 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_input_pipe1_1413_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_input_pipe1_1413_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_input_pipe1_1413_update_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_input_pipe1_1413_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(76), ack => RPIPE_input_pipe1_1413_inst_req_1); -- 
    convolve_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(17) & convolve_CP_3268_elements(77) & convolve_CP_3268_elements(95);
      gj_convolve_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	76 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_input_pipe1_1413_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_input_pipe1_1413_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_input_pipe1_1413_sample_completed_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_input_pipe1_1413_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1413_inst_ack_0, ack => convolve_CP_3268_elements(77)); -- 
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	93 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: 	75 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_input_pipe1_1413_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_input_pipe1_1413_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_input_pipe1_1413_update_completed_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(78) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_input_pipe1_1413_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1413_inst_ack_1, ack => convolve_CP_3268_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	14 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	82 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_kernel_pipe1_1421_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_kernel_pipe1_1421_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_kernel_pipe1_1421_Sample/rr
      -- 
    -- logger for CP element group convolve_CP_3268_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_kernel_pipe1_1421_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(79), ack => RPIPE_kernel_pipe1_1421_inst_req_0); -- 
    convolve_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(14) & convolve_CP_3268_elements(82);
      gj_convolve_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	17 
    -- CP-element group 80: 	81 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	88 
    -- CP-element group 80: 	95 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_kernel_pipe1_1421_update_start_
      -- CP-element group 80: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_kernel_pipe1_1421_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_kernel_pipe1_1421_Update/$entry
      -- 
    -- logger for CP element group convolve_CP_3268_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_kernel_pipe1_1421_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(80), ack => RPIPE_kernel_pipe1_1421_inst_req_1); -- 
    convolve_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(17) & convolve_CP_3268_elements(81) & convolve_CP_3268_elements(88) & convolve_CP_3268_elements(95);
      gj_convolve_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	80 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_kernel_pipe1_1421_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_kernel_pipe1_1421_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_kernel_pipe1_1421_Sample/ra
      -- 
    -- logger for CP element group convolve_CP_3268_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(81) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_kernel_pipe1_1421_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1421_inst_ack_0, ack => convolve_CP_3268_elements(81)); -- 
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	87 
    -- CP-element group 82: 	93 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	37 
    -- CP-element group 82: 	79 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_kernel_pipe1_1421_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_kernel_pipe1_1421_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/RPIPE_kernel_pipe1_1421_Update/$exit
      -- 
    -- logger for CP element group convolve_CP_3268_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:RPIPE_kernel_pipe1_1421_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1421_inst_ack_1, ack => convolve_CP_3268_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	14 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/SUB_u32_u32_1435_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/SUB_u32_u32_1435_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/SUB_u32_u32_1435_sample_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(83) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:SUB_u32_u32_1435_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(83), ack => SUB_u32_u32_1435_inst_req_0); -- 
    convolve_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(14) & convolve_CP_3268_elements(85);
      gj_convolve_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	17 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	91 
    -- CP-element group 84: 	95 
    -- CP-element group 84: 	98 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/SUB_u32_u32_1435_Update/cr
      -- CP-element group 84: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/SUB_u32_u32_1435_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/SUB_u32_u32_1435_update_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(84) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:SUB_u32_u32_1435_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(84), ack => SUB_u32_u32_1435_inst_req_1); -- 
    convolve_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(17) & convolve_CP_3268_elements(91) & convolve_CP_3268_elements(95) & convolve_CP_3268_elements(98);
      gj_convolve_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/SUB_u32_u32_1435_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/SUB_u32_u32_1435_Sample/ra
      -- CP-element group 85: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/SUB_u32_u32_1435_Sample/$exit
      -- 
    -- logger for CP element group convolve_CP_3268_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(85) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:SUB_u32_u32_1435_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_1435_inst_ack_0, ack => convolve_CP_3268_elements(85)); -- 
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	90 
    -- CP-element group 86: 	93 
    -- CP-element group 86: 	97 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	20 
    -- CP-element group 86: 	37 
    -- CP-element group 86: 	56 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/SUB_u32_u32_1435_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/SUB_u32_u32_1435_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/SUB_u32_u32_1435_Update/ca
      -- 
    -- logger for CP element group convolve_CP_3268_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(86) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:SUB_u32_u32_1435_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_1435_inst_ack_1, ack => convolve_CP_3268_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	61 
    -- CP-element group 87: 	82 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	89 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_kernel_pipe1_1469_Sample/req
      -- CP-element group 87: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_kernel_pipe1_1469_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_kernel_pipe1_1469_sample_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(87) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:WPIPE_kernel_pipe1_1469_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(87), ack => WPIPE_kernel_pipe1_1469_inst_req_0); -- 
    convolve_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(61) & convolve_CP_3268_elements(82) & convolve_CP_3268_elements(89);
      gj_convolve_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	57 
    -- CP-element group 88: 	80 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_kernel_pipe1_1469_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_kernel_pipe1_1469_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_kernel_pipe1_1469_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_kernel_pipe1_1469_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_kernel_pipe1_1469_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_kernel_pipe1_1469_Sample/ack
      -- 
    -- logger for CP element group convolve_CP_3268_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:WPIPE_kernel_pipe1_1469_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:WPIPE_kernel_pipe1_1469_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1469_inst_ack_0, ack => convolve_CP_3268_elements(88)); -- 
    req_3517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(88), ack => WPIPE_kernel_pipe1_1469_inst_req_1); -- 
    -- CP-element group 89:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	101 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	87 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_kernel_pipe1_1469_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_kernel_pipe1_1469_Update/ack
      -- CP-element group 89: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_kernel_pipe1_1469_Update/$exit
      -- 
    -- logger for CP element group convolve_CP_3268_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:WPIPE_kernel_pipe1_1469_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1469_inst_ack_1, ack => convolve_CP_3268_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	23 
    -- CP-element group 90: 	61 
    -- CP-element group 90: 	86 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_input_done_pipe_1490_Sample/req
      -- CP-element group 90: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_input_done_pipe_1490_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_input_done_pipe_1490_sample_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(90) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:WPIPE_input_done_pipe_1490_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(90), ack => WPIPE_input_done_pipe_1490_inst_req_0); -- 
    convolve_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(23) & convolve_CP_3268_elements(61) & convolve_CP_3268_elements(86) & convolve_CP_3268_elements(92);
      gj_convolve_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	21 
    -- CP-element group 91: 	57 
    -- CP-element group 91: 	84 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_input_done_pipe_1490_Update/req
      -- CP-element group 91: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_input_done_pipe_1490_update_start_
      -- CP-element group 91: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_input_done_pipe_1490_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_input_done_pipe_1490_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_input_done_pipe_1490_Sample/ack
      -- CP-element group 91: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_input_done_pipe_1490_Sample/$exit
      -- 
    -- logger for CP element group convolve_CP_3268_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(91) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:WPIPE_input_done_pipe_1490_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:WPIPE_input_done_pipe_1490_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1490_inst_ack_0, ack => convolve_CP_3268_elements(91)); -- 
    req_3531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(91), ack => WPIPE_input_done_pipe_1490_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	101 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_input_done_pipe_1490_Update/ack
      -- CP-element group 92: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_input_done_pipe_1490_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_input_done_pipe_1490_Update/$exit
      -- 
    -- logger for CP element group convolve_CP_3268_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(92) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:WPIPE_input_done_pipe_1490_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1490_inst_ack_1, ack => convolve_CP_3268_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	23 
    -- CP-element group 93: 	42 
    -- CP-element group 93: 	78 
    -- CP-element group 93: 	82 
    -- CP-element group 93: 	86 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1496_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1496_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1496_Sample/rr
      -- 
    -- logger for CP element group convolve_CP_3268_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:type_cast_1496_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(93), ack => type_cast_1496_inst_req_0); -- 
    convolve_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(23) & convolve_CP_3268_elements(42) & convolve_CP_3268_elements(78) & convolve_CP_3268_elements(82) & convolve_CP_3268_elements(86) & convolve_CP_3268_elements(95);
      gj_convolve_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	98 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1496_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1496_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1496_update_start_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:type_cast_1496_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(94), ack => type_cast_1496_inst_req_1); -- 
    convolve_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_3268_elements(98);
      gj_convolve_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	21 
    -- CP-element group 95: 	38 
    -- CP-element group 95: 	76 
    -- CP-element group 95: 	80 
    -- CP-element group 95: 	84 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1496_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1496_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1496_Sample/$exit
      -- 
    -- logger for CP element group convolve_CP_3268_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(95) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:type_cast_1496_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1496_inst_ack_0, ack => convolve_CP_3268_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1496_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1496_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/type_cast_1496_update_completed_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(96) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:type_cast_1496_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1496_inst_ack_1, ack => convolve_CP_3268_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	23 
    -- CP-element group 97: 	86 
    -- CP-element group 97: 	96 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_maxpool_output_pipe_1494_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_maxpool_output_pipe_1494_Sample/req
      -- CP-element group 97: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_maxpool_output_pipe_1494_Sample/$entry
      -- 
    -- logger for CP element group convolve_CP_3268_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(97) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:WPIPE_maxpool_output_pipe_1494_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(97), ack => WPIPE_maxpool_output_pipe_1494_inst_req_0); -- 
    convolve_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(23) & convolve_CP_3268_elements(86) & convolve_CP_3268_elements(96) & convolve_CP_3268_elements(99);
      gj_convolve_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	21 
    -- CP-element group 98: 	84 
    -- CP-element group 98: 	94 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_maxpool_output_pipe_1494_Sample/ack
      -- CP-element group 98: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_maxpool_output_pipe_1494_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_maxpool_output_pipe_1494_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_maxpool_output_pipe_1494_update_start_
      -- CP-element group 98: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_maxpool_output_pipe_1494_Update/req
      -- CP-element group 98: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_maxpool_output_pipe_1494_sample_completed_
      -- 
    -- logger for CP element group convolve_CP_3268_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:WPIPE_maxpool_output_pipe_1494_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:WPIPE_maxpool_output_pipe_1494_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1494_inst_ack_0, ack => convolve_CP_3268_elements(98)); -- 
    req_3559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3268_elements(98), ack => WPIPE_maxpool_output_pipe_1494_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_maxpool_output_pipe_1494_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_maxpool_output_pipe_1494_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/WPIPE_maxpool_output_pipe_1494_Update/ack
      -- 
    -- logger for CP element group convolve_CP_3268_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(99) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:WPIPE_maxpool_output_pipe_1494_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1494_inst_ack_1, ack => convolve_CP_3268_elements(99)); -- 
    -- CP-element group 100:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	14 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	15 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group convolve_CP_3268_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(100) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group convolve_CP_3268_elements(100) is a control-delay.
    cp_element_100_delay: control_delay_element  generic map(name => " 100_delay", delay_value => 1)  port map(req => convolve_CP_3268_elements(14), ack => convolve_CP_3268_elements(100), clk => clk, reset =>reset);
    -- CP-element group 101:  join  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	89 
    -- CP-element group 101: 	92 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	11 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1380/do_while_stmt_1396/do_while_stmt_1396_loop_body/$exit
      -- 
    -- logger for CP element group convolve_CP_3268_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(101) fired."); 
        -- 
      end if; --
    end process; 
    convolve_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3268_elements(89) & convolve_CP_3268_elements(92) & convolve_CP_3268_elements(99);
      gj_convolve_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3268_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	10 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1380/do_while_stmt_1396/loop_exit/$exit
      -- CP-element group 102: 	 branch_block_stmt_1380/do_while_stmt_1396/loop_exit/ack
      -- 
    -- logger for CP element group convolve_CP_3268_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(102) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:do_while_stmt_1396_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1396_branch_ack_0, ack => convolve_CP_3268_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	10 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1380/do_while_stmt_1396/loop_taken/$exit
      -- CP-element group 103: 	 branch_block_stmt_1380/do_while_stmt_1396/loop_taken/ack
      -- 
    -- logger for CP element group convolve_CP_3268_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(103) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:do_while_stmt_1396_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1396_branch_ack_1, ack => convolve_CP_3268_elements(103)); -- 
    -- CP-element group 104:  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	8 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	1 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1380/do_while_stmt_1396/$exit
      -- 
    -- logger for CP element group convolve_CP_3268_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and convolve_CP_3268_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:convolve:CP:convolve_CP_3268_elements(104) fired."); 
        -- 
      end if; --
    end process; 
    convolve_CP_3268_elements(104) <= convolve_CP_3268_elements(8);
    convolve_do_while_stmt_1396_terminator_3570: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_1396_terminator_3570", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_3268_elements(11),loop_continue => convolve_CP_3268_elements(103),loop_terminate => convolve_CP_3268_elements(102),loop_back => convolve_CP_3268_elements(9),loop_exit => convolve_CP_3268_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_1398_phi_seq_3374_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_3268_elements(26);
      convolve_CP_3268_elements(29)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_3268_elements(29);
      convolve_CP_3268_elements(30)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_3268_elements(31);
      convolve_CP_3268_elements(27) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_3268_elements(24);
      convolve_CP_3268_elements(33)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_3268_elements(35);
      convolve_CP_3268_elements(34)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_3268_elements(36);
      convolve_CP_3268_elements(25) <= phi_mux_reqs(1);
      phi_stmt_1398_phi_seq_3374 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1398_phi_seq_3374") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_3268_elements(16), 
          phi_sample_ack => convolve_CP_3268_elements(22), 
          phi_update_req => convolve_CP_3268_elements(18), 
          phi_update_ack => convolve_CP_3268_elements(23), 
          phi_mux_ack => convolve_CP_3268_elements(28), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1402_phi_seq_3418_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_3268_elements(45);
      convolve_CP_3268_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_3268_elements(48);
      convolve_CP_3268_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_3268_elements(50);
      convolve_CP_3268_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_3268_elements(43);
      convolve_CP_3268_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_3268_elements(54);
      convolve_CP_3268_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_3268_elements(55);
      convolve_CP_3268_elements(44) <= phi_mux_reqs(1);
      phi_stmt_1402_phi_seq_3418 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1402_phi_seq_3418") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_3268_elements(39), 
          phi_sample_ack => convolve_CP_3268_elements(40), 
          phi_update_req => convolve_CP_3268_elements(41), 
          phi_update_ack => convolve_CP_3268_elements(42), 
          phi_mux_ack => convolve_CP_3268_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1406_phi_seq_3462_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_3268_elements(64);
      convolve_CP_3268_elements(67)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_3268_elements(67);
      convolve_CP_3268_elements(68)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_3268_elements(69);
      convolve_CP_3268_elements(65) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_3268_elements(62);
      convolve_CP_3268_elements(71)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_3268_elements(73);
      convolve_CP_3268_elements(72)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_3268_elements(74);
      convolve_CP_3268_elements(63) <= phi_mux_reqs(1);
      phi_stmt_1406_phi_seq_3462 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1406_phi_seq_3462") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_3268_elements(58), 
          phi_sample_ack => convolve_CP_3268_elements(59), 
          phi_update_req => convolve_CP_3268_elements(60), 
          phi_update_ack => convolve_CP_3268_elements(61), 
          phi_mux_ack => convolve_CP_3268_elements(66), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3326_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_3268_elements(12);
        preds(1)  <= convolve_CP_3268_elements(13);
        entry_tmerge_3326 : transition_merge -- 
          generic map(name => " entry_tmerge_3326")
          port map (preds => preds, symbol_out => convolve_CP_3268_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_1479_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_1460_wire : std_logic_vector(31 downto 0);
    signal MUX_1480_wire : std_logic_vector(15 downto 0);
    signal SUB_u32_u32_1415_1415_delayed_1_0_1436 : std_logic_vector(31 downto 0);
    signal acc_1402 : std_logic_vector(31 downto 0);
    signal acc_val_1448 : std_logic_vector(31 downto 0);
    signal acc_var_1395 : std_logic_vector(31 downto 0);
    signal all_done_flag_1488 : std_logic_vector(0 downto 0);
    signal iread_1414 : std_logic_vector(15 downto 0);
    signal ival_1419 : std_logic_vector(15 downto 0);
    signal konst_1434_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1451_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1457_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1459_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1478_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1491_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1499_wire_constant : std_logic_vector(0 downto 0);
    signal kread_1422 : std_logic_vector(15 downto 0);
    signal kval_1426 : std_logic_vector(15 downto 0);
    signal mcount_var_1390 : std_logic_vector(31 downto 0);
    signal mul_val_1431 : std_logic_vector(15 downto 0);
    signal mycount_1398 : std_logic_vector(31 downto 0);
    signal n_out_count_1483 : std_logic_vector(15 downto 0);
    signal n_out_count_1483_1410_buffered : std_logic_vector(15 downto 0);
    signal nacc_1454 : std_logic_vector(31 downto 0);
    signal nacc_1454_1405_buffered : std_logic_vector(31 downto 0);
    signal next_sum_1441 : std_logic_vector(0 downto 0);
    signal nmycount_1462 : std_logic_vector(31 downto 0);
    signal nmycount_1462_1401_buffered : std_logic_vector(31 downto 0);
    signal num_out_1383 : std_logic_vector(15 downto 0);
    signal out_count_1406 : std_logic_vector(15 downto 0);
    signal out_done_flag_1467 : std_logic_vector(0 downto 0);
    signal size_1386 : std_logic_vector(31 downto 0);
    signal type_cast_1409_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1444_wire : std_logic_vector(31 downto 0);
    signal type_cast_1446_wire : std_logic_vector(31 downto 0);
    signal type_cast_1476_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1496_wire : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    acc_var_1395 <= "00000000000000000000000000000000";
    konst_1434_wire_constant <= "00000000000000000000000000000001";
    konst_1451_wire_constant <= "00000000000000000000000000000000";
    konst_1457_wire_constant <= "00000000000000000000000000000000";
    konst_1459_wire_constant <= "00000000000000000000000000000001";
    konst_1478_wire_constant <= "0000000000000001";
    konst_1491_wire_constant <= "1";
    konst_1499_wire_constant <= "1";
    mcount_var_1390 <= "00000000000000000000000000000000";
    type_cast_1409_wire_constant <= "0000000000000001";
    type_cast_1476_wire_constant <= "0000000000000001";
    -- logger for phi phi_stmt_1398
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1398_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolve:DP:phi_stmt_1398:input-0 mcount_var_1390= " & Convert_SLV_To_Hex_String(mcount_var_1390));
          --
        end if;
        if phi_stmt_1398_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolve:DP:phi_stmt_1398:input-1 nmycount_1462_1401_buffered= " & Convert_SLV_To_Hex_String(nmycount_1462_1401_buffered));
          --
        end if;
        if phi_stmt_1398_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolve:DP:phi_stmt_1398:sample-completed");
          --
        end if;
        if phi_stmt_1398_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolve:DP:phi_stmt_1398:output mycount_1398= " & Convert_SLV_To_Hex_String(mycount_1398));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1398: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= mcount_var_1390 & nmycount_1462_1401_buffered;
      req <= phi_stmt_1398_req_0 & phi_stmt_1398_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1398",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1398_ack_0,
          idata => idata,
          odata => mycount_1398,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1398
    -- logger for phi phi_stmt_1402
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1402_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolve:DP:phi_stmt_1402:input-0 acc_var_1395= " & Convert_SLV_To_Hex_String(acc_var_1395));
          --
        end if;
        if phi_stmt_1402_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolve:DP:phi_stmt_1402:input-1 nacc_1454_1405_buffered= " & Convert_SLV_To_Hex_String(nacc_1454_1405_buffered));
          --
        end if;
        if phi_stmt_1402_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolve:DP:phi_stmt_1402:sample-completed");
          --
        end if;
        if phi_stmt_1402_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolve:DP:phi_stmt_1402:output acc_1402= " & Convert_SLV_To_Hex_String(acc_1402));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1402: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= acc_var_1395 & nacc_1454_1405_buffered;
      req <= phi_stmt_1402_req_0 & phi_stmt_1402_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1402",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1402_ack_0,
          idata => idata,
          odata => acc_1402,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1402
    -- logger for phi phi_stmt_1406
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1406_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolve:DP:phi_stmt_1406:input-0 type_cast_1409_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1409_wire_constant));
          --
        end if;
        if phi_stmt_1406_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:convolve:DP:phi_stmt_1406:input-1 n_out_count_1483_1410_buffered= " & Convert_SLV_To_Hex_String(n_out_count_1483_1410_buffered));
          --
        end if;
        if phi_stmt_1406_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:convolve:DP:phi_stmt_1406:sample-completed");
          --
        end if;
        if phi_stmt_1406_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:convolve:DP:phi_stmt_1406:output out_count_1406= " & Convert_SLV_To_Hex_String(out_count_1406));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1406: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1409_wire_constant & n_out_count_1483_1410_buffered;
      req <= phi_stmt_1406_req_0 & phi_stmt_1406_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1406",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1406_ack_0,
          idata => idata,
          odata => out_count_1406,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1406
    -- logger for split-operator MUX_1453_inst flow-through 
    process(nacc_1454) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:MUX_1453_inst:flowthrough inputs: " & " next_sum_1441 = "& Convert_SLV_To_Hex_String(next_sum_1441) & " konst_1451_wire_constant = "& Convert_SLV_To_Hex_String(konst_1451_wire_constant) & " acc_val_1448 = "& Convert_SLV_To_Hex_String(acc_val_1448) & " outputs:" & " nacc_1454= "  & Convert_SLV_To_Hex_String(nacc_1454));
      --
    end process; 
    -- flow-through select operator MUX_1453_inst
    nacc_1454 <= konst_1451_wire_constant when (next_sum_1441(0) /=  '0') else acc_val_1448;
    -- logger for split-operator MUX_1461_inst flow-through 
    process(nmycount_1462) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:MUX_1461_inst:flowthrough inputs: " & " next_sum_1441 = "& Convert_SLV_To_Hex_String(next_sum_1441) & " konst_1457_wire_constant = "& Convert_SLV_To_Hex_String(konst_1457_wire_constant) & " ADD_u32_u32_1460_wire = "& Convert_SLV_To_Hex_String(ADD_u32_u32_1460_wire) & " outputs:" & " nmycount_1462= "  & Convert_SLV_To_Hex_String(nmycount_1462));
      --
    end process; 
    -- flow-through select operator MUX_1461_inst
    nmycount_1462 <= konst_1457_wire_constant when (next_sum_1441(0) /=  '0') else ADD_u32_u32_1460_wire;
    -- logger for split-operator MUX_1480_inst flow-through 
    process(MUX_1480_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:MUX_1480_inst:flowthrough inputs: " & " out_done_flag_1467 = "& Convert_SLV_To_Hex_String(out_done_flag_1467) & " type_cast_1476_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1476_wire_constant) & " ADD_u16_u16_1479_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1479_wire) & " outputs:" & " MUX_1480_wire= "  & Convert_SLV_To_Hex_String(MUX_1480_wire));
      --
    end process; 
    -- flow-through select operator MUX_1480_inst
    MUX_1480_wire <= type_cast_1476_wire_constant when (out_done_flag_1467(0) /=  '0') else ADD_u16_u16_1479_wire;
    -- logger for split-operator MUX_1482_inst flow-through 
    process(n_out_count_1483) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:MUX_1482_inst:flowthrough inputs: " & " next_sum_1441 = "& Convert_SLV_To_Hex_String(next_sum_1441) & " MUX_1480_wire = "& Convert_SLV_To_Hex_String(MUX_1480_wire) & " out_count_1406 = "& Convert_SLV_To_Hex_String(out_count_1406) & " outputs:" & " n_out_count_1483= "  & Convert_SLV_To_Hex_String(n_out_count_1483));
      --
    end process; 
    -- flow-through select operator MUX_1482_inst
    n_out_count_1483 <= MUX_1480_wire when (next_sum_1441(0) /=  '0') else out_count_1406;
    -- logger for split-operator n_out_count_1483_1410_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_out_count_1483_1410_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:n_out_count_1483_1410_buf:started:   inputs: " & " n_out_count_1483 = "& Convert_SLV_To_Hex_String(n_out_count_1483));
          --
        end if; 
        if n_out_count_1483_1410_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:n_out_count_1483_1410_buf:finished:  outputs: " & " n_out_count_1483_1410_buffered= "  & Convert_SLV_To_Hex_String(n_out_count_1483_1410_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_out_count_1483_1410_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_out_count_1483_1410_buf_req_0;
      n_out_count_1483_1410_buf_ack_0<= wack(0);
      rreq(0) <= n_out_count_1483_1410_buf_req_1;
      n_out_count_1483_1410_buf_ack_1<= rack(0);
      n_out_count_1483_1410_buf : InterlockBuffer generic map ( -- 
        name => "n_out_count_1483_1410_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_out_count_1483,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_out_count_1483_1410_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator nacc_1454_1405_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if nacc_1454_1405_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:nacc_1454_1405_buf:started:   inputs: " & " nacc_1454 = "& Convert_SLV_To_Hex_String(nacc_1454));
          --
        end if; 
        if nacc_1454_1405_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:nacc_1454_1405_buf:finished:  outputs: " & " nacc_1454_1405_buffered= "  & Convert_SLV_To_Hex_String(nacc_1454_1405_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    nacc_1454_1405_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc_1454_1405_buf_req_0;
      nacc_1454_1405_buf_ack_0<= wack(0);
      rreq(0) <= nacc_1454_1405_buf_req_1;
      nacc_1454_1405_buf_ack_1<= rack(0);
      nacc_1454_1405_buf : InterlockBuffer generic map ( -- 
        name => "nacc_1454_1405_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc_1454,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc_1454_1405_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator nmycount_1462_1401_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if nmycount_1462_1401_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:nmycount_1462_1401_buf:started:   inputs: " & " nmycount_1462 = "& Convert_SLV_To_Hex_String(nmycount_1462));
          --
        end if; 
        if nmycount_1462_1401_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:nmycount_1462_1401_buf:finished:  outputs: " & " nmycount_1462_1401_buffered= "  & Convert_SLV_To_Hex_String(nmycount_1462_1401_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    nmycount_1462_1401_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_1462_1401_buf_req_0;
      nmycount_1462_1401_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_1462_1401_buf_req_1;
      nmycount_1462_1401_buf_ack_1<= rack(0);
      nmycount_1462_1401_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_1462_1401_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_1462,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_1462_1401_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1418_inst flow-through 
    process(ival_1419) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:type_cast_1418_inst:flowthrough inputs: " & " iread_1414 = "& Convert_SLV_To_Hex_String(iread_1414) & " outputs:" & " ival_1419= "  & Convert_SLV_To_Hex_String(ival_1419));
      --
    end process; 
    -- interlock type_cast_1418_inst
    process(iread_1414) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread_1414(15 downto 0);
      ival_1419 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1425_inst flow-through 
    process(kval_1426) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:type_cast_1425_inst:flowthrough inputs: " & " kread_1422 = "& Convert_SLV_To_Hex_String(kread_1422) & " outputs:" & " kval_1426= "  & Convert_SLV_To_Hex_String(kval_1426));
      --
    end process; 
    -- interlock type_cast_1425_inst
    process(kread_1422) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread_1422(15 downto 0);
      kval_1426 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1444_inst flow-through 
    process(type_cast_1444_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:type_cast_1444_inst:flowthrough inputs: " & " acc_1402 = "& Convert_SLV_To_Hex_String(acc_1402) & " outputs:" & " type_cast_1444_wire= "  & Convert_SLV_To_Hex_String(type_cast_1444_wire));
      --
    end process; 
    -- interlock type_cast_1444_inst
    process(acc_1402) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := acc_1402(31 downto 0);
      type_cast_1444_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1446_inst flow-through 
    process(type_cast_1446_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:type_cast_1446_inst:flowthrough inputs: " & " mul_val_1431 = "& Convert_SLV_To_Hex_String(mul_val_1431) & " outputs:" & " type_cast_1446_wire= "  & Convert_SLV_To_Hex_String(type_cast_1446_wire));
      --
    end process; 
    -- interlock type_cast_1446_inst
    process(mul_val_1431) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := mul_val_1431(15 downto 0);
      type_cast_1446_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1496_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1496_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:type_cast_1496_inst:started:   inputs: " & " next_sum_1441 (guard)= " & Convert_SLV_To_String(next_sum_1441) & " acc_val_1448 = "& Convert_SLV_To_Hex_String(acc_val_1448));
          --
        end if; 
        if type_cast_1496_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:type_cast_1496_inst:finished:  outputs: " & " type_cast_1496_wire= "  & Convert_SLV_To_Hex_String(type_cast_1496_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1496_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1496_inst_req_0;
      type_cast_1496_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1496_inst_req_1;
      type_cast_1496_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1441(0);
      type_cast_1496_inst_gI: SplitGuardInterface generic map(name => "type_cast_1496_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1496_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1496_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_1448,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1496_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1396_branch_req_0," req0 do_while_stmt_1396_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1396_branch_ack_0," ack0 do_while_stmt_1396_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1396_branch_ack_1," ack1 do_while_stmt_1396_branch");
    do_while_stmt_1396_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1499_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1396_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1396_branch_req_0,
          ack0 => do_while_stmt_1396_branch_ack_0,
          ack1 => do_while_stmt_1396_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_i32_i32_1447_inst flow-through 
    process(acc_val_1448) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:ADD_i32_i32_1447_inst:flowthrough inputs: " & " type_cast_1444_wire = "& Convert_SLV_To_Hex_String(type_cast_1444_wire) & " type_cast_1446_wire = "& Convert_SLV_To_Hex_String(type_cast_1446_wire) & " outputs:" & " acc_val_1448= "  & Convert_SLV_To_Hex_String(acc_val_1448));
      --
    end process; 
    -- binary operator ADD_i32_i32_1447_inst
    process(type_cast_1444_wire, type_cast_1446_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(type_cast_1444_wire, type_cast_1446_wire, tmp_var);
      acc_val_1448 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1479_inst flow-through 
    process(ADD_u16_u16_1479_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:ADD_u16_u16_1479_inst:flowthrough inputs: " & " out_count_1406 = "& Convert_SLV_To_Hex_String(out_count_1406) & " konst_1478_wire_constant = "& Convert_SLV_To_Hex_String(konst_1478_wire_constant) & " outputs:" & " ADD_u16_u16_1479_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1479_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1479_inst
    process(out_count_1406) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(out_count_1406, konst_1478_wire_constant, tmp_var);
      ADD_u16_u16_1479_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1460_inst flow-through 
    process(ADD_u32_u32_1460_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:ADD_u32_u32_1460_inst:flowthrough inputs: " & " mycount_1398 = "& Convert_SLV_To_Hex_String(mycount_1398) & " konst_1459_wire_constant = "& Convert_SLV_To_Hex_String(konst_1459_wire_constant) & " outputs:" & " ADD_u32_u32_1460_wire= "  & Convert_SLV_To_Hex_String(ADD_u32_u32_1460_wire));
      --
    end process; 
    -- binary operator ADD_u32_u32_1460_inst
    process(mycount_1398) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_1398, konst_1459_wire_constant, tmp_var);
      ADD_u32_u32_1460_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_1487_inst flow-through 
    process(all_done_flag_1488) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:AND_u1_u1_1487_inst:flowthrough inputs: " & " out_done_flag_1467 = "& Convert_SLV_To_Hex_String(out_done_flag_1467) & " next_sum_1441 = "& Convert_SLV_To_Hex_String(next_sum_1441) & " outputs:" & " all_done_flag_1488= "  & Convert_SLV_To_Hex_String(all_done_flag_1488));
      --
    end process; 
    -- binary operator AND_u1_u1_1487_inst
    process(out_done_flag_1467, next_sum_1441) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_1467, next_sum_1441, tmp_var);
      all_done_flag_1488 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u16_u1_1466_inst flow-through 
    process(out_done_flag_1467) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:EQ_u16_u1_1466_inst:flowthrough inputs: " & " out_count_1406 = "& Convert_SLV_To_Hex_String(out_count_1406) & " num_out_1383 = "& Convert_SLV_To_Hex_String(num_out_1383) & " outputs:" & " out_done_flag_1467= "  & Convert_SLV_To_Hex_String(out_done_flag_1467));
      --
    end process; 
    -- binary operator EQ_u16_u1_1466_inst
    process(out_count_1406, num_out_1383) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(out_count_1406, num_out_1383, tmp_var);
      out_done_flag_1467 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u32_u1_1440_inst flow-through 
    process(next_sum_1441) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:EQ_u32_u1_1440_inst:flowthrough inputs: " & " mycount_1398 = "& Convert_SLV_To_Hex_String(mycount_1398) & " SUB_u32_u32_1415_1415_delayed_1_0_1436 = "& Convert_SLV_To_Hex_String(SUB_u32_u32_1415_1415_delayed_1_0_1436) & " outputs:" & " next_sum_1441= "  & Convert_SLV_To_Hex_String(next_sum_1441));
      --
    end process; 
    -- binary operator EQ_u32_u1_1440_inst
    process(mycount_1398, SUB_u32_u32_1415_1415_delayed_1_0_1436) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycount_1398, SUB_u32_u32_1415_1415_delayed_1_0_1436, tmp_var);
      next_sum_1441 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_i16_i16_1430_inst flow-through 
    process(mul_val_1431) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:MUL_i16_i16_1430_inst:flowthrough inputs: " & " kval_1426 = "& Convert_SLV_To_Hex_String(kval_1426) & " ival_1419 = "& Convert_SLV_To_Hex_String(ival_1419) & " outputs:" & " mul_val_1431= "  & Convert_SLV_To_Hex_String(mul_val_1431));
      --
    end process; 
    -- binary operator MUL_i16_i16_1430_inst
    process(kval_1426, ival_1419) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval_1426, ival_1419, tmp_var);
      mul_val_1431 <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u32_u32_1435_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if SUB_u32_u32_1435_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:SUB_u32_u32_1435_inst:started:   inputs: " & " size_1386 = "& Convert_SLV_To_Hex_String(size_1386) & " konst_1434_wire_constant = "& Convert_SLV_To_Hex_String(konst_1434_wire_constant));
          --
        end if; 
        if SUB_u32_u32_1435_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:SUB_u32_u32_1435_inst:finished:  outputs: " & " SUB_u32_u32_1415_1415_delayed_1_0_1436= "  & Convert_SLV_To_Hex_String(SUB_u32_u32_1415_1415_delayed_1_0_1436));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (7) : SUB_u32_u32_1435_inst 
    ApIntSub_group_7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= size_1386;
      SUB_u32_u32_1415_1415_delayed_1_0_1436 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_1435_inst_req_0;
      SUB_u32_u32_1435_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_1435_inst_req_1;
      SUB_u32_u32_1435_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_7_gI: SplitGuardInterface generic map(name => "ApIntSub_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- logger for split-operator RPIPE_input_pipe1_1413_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_input_pipe1_1413_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:RPIPE_input_pipe1_1413_inst:started:   PipeRead from input_pipe1 inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_input_pipe1_1413_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:RPIPE_input_pipe1_1413_inst:finished:  outputs: " & " iread_1414= "  & Convert_SLV_To_Hex_String(iread_1414));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_input_pipe1_1413_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_1413_inst_req_0;
      RPIPE_input_pipe1_1413_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_1413_inst_req_1;
      RPIPE_input_pipe1_1413_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iread_1414 <= data_out(15 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator RPIPE_kernel_pipe1_1421_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_kernel_pipe1_1421_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:RPIPE_kernel_pipe1_1421_inst:started:   PipeRead from kernel_pipe1 inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_kernel_pipe1_1421_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:RPIPE_kernel_pipe1_1421_inst:finished:  outputs: " & " kread_1422= "  & Convert_SLV_To_Hex_String(kread_1422));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (1) : RPIPE_kernel_pipe1_1421_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_1421_inst_req_0;
      RPIPE_kernel_pipe1_1421_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_1421_inst_req_1;
      RPIPE_kernel_pipe1_1421_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      kread_1422 <= data_out(15 downto 0);
      kernel_pipe1_read_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_1: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- logger for split-operator RPIPE_num_out_pipe_1382_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_num_out_pipe_1382_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:RPIPE_num_out_pipe_1382_inst:started:   PipeRead from num_out_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_num_out_pipe_1382_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:RPIPE_num_out_pipe_1382_inst:finished:  outputs: " & " num_out_1383= "  & Convert_SLV_To_Hex_String(num_out_1383));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (2) : RPIPE_num_out_pipe_1382_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_num_out_pipe_1382_inst_req_0;
      RPIPE_num_out_pipe_1382_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_num_out_pipe_1382_inst_req_1;
      RPIPE_num_out_pipe_1382_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      num_out_1383 <= data_out(15 downto 0);
      num_out_pipe_read_2_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_2: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- logger for split-operator RPIPE_size_pipe_1385_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_size_pipe_1385_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:RPIPE_size_pipe_1385_inst:started:   PipeRead from size_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_size_pipe_1385_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:RPIPE_size_pipe_1385_inst:finished:  outputs: " & " size_1386= "  & Convert_SLV_To_Hex_String(size_1386));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (3) : RPIPE_size_pipe_1385_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_1385_inst_req_0;
      RPIPE_size_pipe_1385_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_1385_inst_req_1;
      RPIPE_size_pipe_1385_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      size_1386 <= data_out(31 downto 0);
      size_pipe_read_3_gI: SplitGuardInterface generic map(name => "size_pipe_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_3: InputPortRevised -- 
        generic map ( name => "size_pipe_read_3", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- logger for split-operator WPIPE_input_done_pipe_1490_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_input_done_pipe_1490_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:WPIPE_input_done_pipe_1490_inst:started:   PipeWrite to input_done_pipe inputs: " & " all_done_flag_1488 (guard)= " & Convert_SLV_To_String(all_done_flag_1488) & " konst_1491_wire_constant = "& Convert_SLV_To_Hex_String(konst_1491_wire_constant));
          --
        end if; 
        if WPIPE_input_done_pipe_1490_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:WPIPE_input_done_pipe_1490_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_input_done_pipe_1490_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_1490_inst_req_0;
      WPIPE_input_done_pipe_1490_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_1490_inst_req_1;
      WPIPE_input_done_pipe_1490_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= all_done_flag_1488(0);
      data_in <= konst_1491_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator WPIPE_kernel_pipe1_1469_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_kernel_pipe1_1469_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:WPIPE_kernel_pipe1_1469_inst:started:   PipeWrite to kernel_pipe1 inputs: " & " out_done_flag_1467 (guard complement )= " & Convert_SLV_To_String(out_done_flag_1467) & " kread_1422 = "& Convert_SLV_To_Hex_String(kread_1422));
          --
        end if; 
        if WPIPE_kernel_pipe1_1469_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:WPIPE_kernel_pipe1_1469_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (1) : WPIPE_kernel_pipe1_1469_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_1469_inst_req_0;
      WPIPE_kernel_pipe1_1469_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_1469_inst_req_1;
      WPIPE_kernel_pipe1_1469_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  not out_done_flag_1467(0);
      data_in <= kread_1422;
      kernel_pipe1_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logger for split-operator WPIPE_maxpool_output_pipe_1494_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_maxpool_output_pipe_1494_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:WPIPE_maxpool_output_pipe_1494_inst:started:   PipeWrite to maxpool_output_pipe inputs: " & " next_sum_1441 (guard)= " & Convert_SLV_To_String(next_sum_1441) & " type_cast_1496_wire = "& Convert_SLV_To_Hex_String(type_cast_1496_wire));
          --
        end if; 
        if WPIPE_maxpool_output_pipe_1494_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:convolve:DP:WPIPE_maxpool_output_pipe_1494_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (2) : WPIPE_maxpool_output_pipe_1494_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1494_inst_req_0;
      WPIPE_maxpool_output_pipe_1494_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1494_inst_req_1;
      WPIPE_maxpool_output_pipe_1494_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= next_sum_1441(0);
      data_in <= type_cast_1496_wire;
      maxpool_output_pipe_write_2_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(63 downto 0);
    end_add : in  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 128)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(63 downto 0);
  signal start_add_update_enable: Boolean;
  signal end_add_buffer :  std_logic_vector(63 downto 0);
  signal end_add_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_676_start: Boolean;
  signal loadKernelChannel_CP_676_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal nfetch_val_418_357_buf_ack_1 : boolean;
  signal array_obj_ref_396_index_offset_req_1 : boolean;
  signal W_fetch_val_395_delayed_13_0_410_inst_ack_0 : boolean;
  signal W_fetch_val_395_delayed_13_0_410_inst_ack_1 : boolean;
  signal array_obj_ref_396_index_offset_ack_1 : boolean;
  signal phi_stmt_355_req_1 : boolean;
  signal W_fn_393_delayed_13_0_407_inst_ack_1 : boolean;
  signal do_while_stmt_349_branch_ack_1 : boolean;
  signal ptr_deref_405_load_0_ack_1 : boolean;
  signal do_while_stmt_349_branch_ack_0 : boolean;
  signal WPIPE_size_pipe_427_inst_req_0 : boolean;
  signal WPIPE_size_pipe_427_inst_req_1 : boolean;
  signal start_add_354_buf_ack_1 : boolean;
  signal start_add_354_buf_req_1 : boolean;
  signal WPIPE_size_pipe_427_inst_ack_1 : boolean;
  signal my_fetch_338_358_buf_req_1 : boolean;
  signal nfetch_val_418_357_buf_ack_0 : boolean;
  signal phi_stmt_355_req_0 : boolean;
  signal my_fetch_338_358_buf_req_0 : boolean;
  signal W_fetch_val_395_delayed_13_0_410_inst_req_1 : boolean;
  signal W_fetch_val_395_delayed_13_0_410_inst_req_0 : boolean;
  signal W_fn_387_delayed_7_0_399_inst_req_0 : boolean;
  signal type_cast_431_inst_req_0 : boolean;
  signal addr_of_397_final_reg_req_0 : boolean;
  signal addr_of_397_final_reg_ack_0 : boolean;
  signal my_fetch_338_358_buf_ack_1 : boolean;
  signal W_fn_393_delayed_13_0_407_inst_req_1 : boolean;
  signal addr_of_397_final_reg_req_1 : boolean;
  signal addr_of_397_final_reg_ack_1 : boolean;
  signal type_cast_431_inst_req_1 : boolean;
  signal phi_stmt_355_ack_0 : boolean;
  signal W_fn_387_delayed_7_0_399_inst_ack_0 : boolean;
  signal nfetch_val_418_357_buf_req_0 : boolean;
  signal W_fn_393_delayed_13_0_407_inst_ack_0 : boolean;
  signal my_fetch_338_358_buf_ack_0 : boolean;
  signal array_obj_ref_396_index_offset_req_0 : boolean;
  signal array_obj_ref_396_index_offset_ack_0 : boolean;
  signal nfetch_val_418_357_buf_req_1 : boolean;
  signal type_cast_431_inst_ack_1 : boolean;
  signal type_cast_431_inst_ack_0 : boolean;
  signal W_fn_393_delayed_13_0_407_inst_req_0 : boolean;
  signal start_add_354_buf_ack_0 : boolean;
  signal ptr_deref_405_load_0_req_1 : boolean;
  signal WPIPE_kernel_pipe1_380_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_380_inst_req_1 : boolean;
  signal start_add_354_buf_req_0 : boolean;
  signal array_obj_ref_332_index_offset_req_0 : boolean;
  signal array_obj_ref_332_index_offset_ack_0 : boolean;
  signal array_obj_ref_332_index_offset_req_1 : boolean;
  signal array_obj_ref_332_index_offset_ack_1 : boolean;
  signal WPIPE_size_pipe_427_inst_ack_0 : boolean;
  signal addr_of_333_final_reg_req_0 : boolean;
  signal addr_of_333_final_reg_ack_0 : boolean;
  signal addr_of_333_final_reg_req_1 : boolean;
  signal addr_of_333_final_reg_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_380_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_380_inst_req_0 : boolean;
  signal ptr_deref_405_load_0_ack_0 : boolean;
  signal ptr_deref_405_load_0_req_0 : boolean;
  signal W_fn_387_delayed_7_0_399_inst_ack_1 : boolean;
  signal W_fn_387_delayed_7_0_399_inst_req_1 : boolean;
  signal ptr_deref_337_load_0_req_0 : boolean;
  signal ptr_deref_337_load_0_ack_0 : boolean;
  signal ptr_deref_337_load_0_req_1 : boolean;
  signal ptr_deref_337_load_0_ack_1 : boolean;
  signal RPIPE_input_done_pipe_346_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_346_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_346_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_346_inst_ack_1 : boolean;
  signal do_while_stmt_349_branch_req_0 : boolean;
  signal phi_stmt_351_req_0 : boolean;
  signal phi_stmt_351_req_1 : boolean;
  signal phi_stmt_351_ack_0 : boolean;
  signal nmycount_373_353_buf_req_0 : boolean;
  signal nmycount_373_353_buf_ack_0 : boolean;
  signal nmycount_373_353_buf_req_1 : boolean;
  signal nmycount_373_353_buf_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 128) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(127 downto 64) <= end_add;
  end_add_buffer <= in_buffer_data_out(127 downto 64);
  in_buffer_data_in(tag_length + 127 downto 128) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 127 downto 128);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_676_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,loadKernelChannel_CP_676_start,"loadKernelChannel cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,loadKernelChannel_CP_676_symbol, "loadKernelChannel cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_676: Block -- control-path 
    signal loadKernelChannel_CP_676_elements: BooleanArray(94 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_676_elements(0) <= loadKernelChannel_CP_676_start;
    loadKernelChannel_CP_676_symbol <= loadKernelChannel_CP_676_elements(94);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/$entry
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/addr_of_333_update_start_
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_index_resized_1
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_index_computed_1
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/addr_of_333_complete/$entry
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/addr_of_333_complete/req
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_update_start_
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Update/$entry
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/RPIPE_input_done_pipe_346_sample_start_
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/RPIPE_input_done_pipe_346_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_327_to_assign_stmt_347/RPIPE_input_done_pipe_346_Sample/rr
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:addr_of_333_final_reg_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:RPIPE_input_done_pipe_346_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:array_obj_ref_332_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:array_obj_ref_332_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:ptr_deref_337_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => addr_of_333_final_reg_req_1); -- 
    rr_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => RPIPE_input_done_pipe_346_inst_req_0); -- 
    req_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => array_obj_ref_332_index_offset_req_0); -- 
    req_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => array_obj_ref_332_index_offset_req_1); -- 
    cr_771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => ptr_deref_337_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_final_index_sum_regn_sample_complete
      -- CP-element group 1: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_final_index_sum_regn_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:array_obj_ref_332_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_332_index_offset_ack_0, ack => loadKernelChannel_CP_676_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_327_to_assign_stmt_347/addr_of_333_sample_start_
      -- CP-element group 2: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_root_address_calculated
      -- CP-element group 2: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_offset_calculated
      -- CP-element group 2: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_final_index_sum_regn_Update/$exit
      -- CP-element group 2: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_final_index_sum_regn_Update/ack
      -- CP-element group 2: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_base_plus_offset/$entry
      -- CP-element group 2: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_base_plus_offset/$exit
      -- CP-element group 2: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 assign_stmt_327_to_assign_stmt_347/array_obj_ref_332_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 assign_stmt_327_to_assign_stmt_347/addr_of_333_request/$entry
      -- CP-element group 2: 	 assign_stmt_327_to_assign_stmt_347/addr_of_333_request/req
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:array_obj_ref_332_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:addr_of_333_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_332_index_offset_ack_1, ack => loadKernelChannel_CP_676_elements(2)); -- 
    req_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(2), ack => addr_of_333_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_327_to_assign_stmt_347/addr_of_333_sample_completed_
      -- CP-element group 3: 	 assign_stmt_327_to_assign_stmt_347/addr_of_333_request/$exit
      -- CP-element group 3: 	 assign_stmt_327_to_assign_stmt_347/addr_of_333_request/ack
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:addr_of_333_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_333_final_reg_ack_0, ack => loadKernelChannel_CP_676_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (24) 
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/addr_of_333_update_completed_
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/addr_of_333_complete/$exit
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/addr_of_333_complete/ack
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_sample_start_
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_base_address_calculated
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_word_address_calculated
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_root_address_calculated
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_base_address_resized
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_base_addr_resize/$entry
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_base_addr_resize/$exit
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_base_plus_offset/$entry
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_base_plus_offset/$exit
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_word_addrgen/$entry
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_word_addrgen/$exit
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_word_addrgen/root_register_req
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_word_addrgen/root_register_ack
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Sample/word_access_start/$entry
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Sample/word_access_start/word_0/$entry
      -- CP-element group 4: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:addr_of_333_final_reg_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:ptr_deref_337_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_333_final_reg_ack_1, ack => loadKernelChannel_CP_676_elements(4)); -- 
    rr_760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(4), ack => ptr_deref_337_load_0_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_sample_completed_
      -- CP-element group 5: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Sample/word_access_start/$exit
      -- CP-element group 5: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:ptr_deref_337_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_337_load_0_ack_0, ack => loadKernelChannel_CP_676_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_update_completed_
      -- CP-element group 6: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Update/$exit
      -- CP-element group 6: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Update/word_access_complete/$exit
      -- CP-element group 6: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Update/ptr_deref_337_Merge/$entry
      -- CP-element group 6: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Update/ptr_deref_337_Merge/$exit
      -- CP-element group 6: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Update/ptr_deref_337_Merge/merge_req
      -- CP-element group 6: 	 assign_stmt_327_to_assign_stmt_347/ptr_deref_337_Update/ptr_deref_337_Merge/merge_ack
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:ptr_deref_337_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_337_load_0_ack_1, ack => loadKernelChannel_CP_676_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_327_to_assign_stmt_347/RPIPE_input_done_pipe_346_sample_completed_
      -- CP-element group 7: 	 assign_stmt_327_to_assign_stmt_347/RPIPE_input_done_pipe_346_update_start_
      -- CP-element group 7: 	 assign_stmt_327_to_assign_stmt_347/RPIPE_input_done_pipe_346_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_327_to_assign_stmt_347/RPIPE_input_done_pipe_346_Sample/ra
      -- CP-element group 7: 	 assign_stmt_327_to_assign_stmt_347/RPIPE_input_done_pipe_346_Update/$entry
      -- CP-element group 7: 	 assign_stmt_327_to_assign_stmt_347/RPIPE_input_done_pipe_346_Update/cr
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:RPIPE_input_done_pipe_346_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:RPIPE_input_done_pipe_346_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_346_inst_ack_0, ack => loadKernelChannel_CP_676_elements(7)); -- 
    cr_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(7), ack => RPIPE_input_done_pipe_346_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_327_to_assign_stmt_347/RPIPE_input_done_pipe_346_update_completed_
      -- CP-element group 8: 	 assign_stmt_327_to_assign_stmt_347/RPIPE_input_done_pipe_346_Update/$exit
      -- CP-element group 8: 	 assign_stmt_327_to_assign_stmt_347/RPIPE_input_done_pipe_346_Update/ca
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:RPIPE_input_done_pipe_346_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_346_inst_ack_1, ack => loadKernelChannel_CP_676_elements(8)); -- 
    -- CP-element group 9:  join  transition  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: 	8 
    -- CP-element group 9: 	1 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 assign_stmt_327_to_assign_stmt_347/$exit
      -- CP-element group 9: 	 branch_block_stmt_348/$entry
      -- CP-element group 9: 	 branch_block_stmt_348/branch_block_stmt_348__entry__
      -- CP-element group 9: 	 branch_block_stmt_348/do_while_stmt_349__entry__
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "loadKernelChannel_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(6) & loadKernelChannel_CP_676_elements(8) & loadKernelChannel_CP_676_elements(1);
      gj_loadKernelChannel_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  place  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	90 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	91 
    -- CP-element group 10: 	92 
    -- CP-element group 10:  members (10) 
      -- CP-element group 10: 	 assign_stmt_432/$entry
      -- CP-element group 10: 	 assign_stmt_432/type_cast_431_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_432/type_cast_431_update_start_
      -- CP-element group 10: 	 assign_stmt_432/type_cast_431_Sample/rr
      -- CP-element group 10: 	 assign_stmt_432/type_cast_431_Update/cr
      -- CP-element group 10: 	 assign_stmt_432/type_cast_431_sample_start_
      -- CP-element group 10: 	 assign_stmt_432/type_cast_431_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_348/$exit
      -- CP-element group 10: 	 branch_block_stmt_348/branch_block_stmt_348__exit__
      -- CP-element group 10: 	 branch_block_stmt_348/do_while_stmt_349__exit__
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:type_cast_431_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:type_cast_431_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    rr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(10), ack => type_cast_431_inst_req_0); -- 
    cr_1104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(10), ack => type_cast_431_inst_req_1); -- 
    loadKernelChannel_CP_676_elements(10) <= loadKernelChannel_CP_676_elements(90);
    -- CP-element group 11:  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_348/do_while_stmt_349/$entry
      -- CP-element group 11: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349__entry__
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_CP_676_elements(11) <= loadKernelChannel_CP_676_elements(9);
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	90 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349__exit__
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group loadKernelChannel_CP_676_elements(12) is bound as output of CP function.
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_348/do_while_stmt_349/loop_back
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group loadKernelChannel_CP_676_elements(13) is bound as output of CP function.
    -- CP-element group 14:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	89 
    -- CP-element group 14: 	88 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_348/do_while_stmt_349/loop_exit/$entry
      -- CP-element group 14: 	 branch_block_stmt_348/do_while_stmt_349/loop_taken/$entry
      -- CP-element group 14: 	 branch_block_stmt_348/do_while_stmt_349/condition_done
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_CP_676_elements(14) <= loadKernelChannel_CP_676_elements(19);
    -- CP-element group 15:  branch  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	87 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_348/do_while_stmt_349/loop_body_done
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_CP_676_elements(15) <= loadKernelChannel_CP_676_elements(87);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	47 
    -- CP-element group 16: 	30 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_CP_676_elements(16) <= loadKernelChannel_CP_676_elements(13);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	49 
    -- CP-element group 17: 	32 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_CP_676_elements(17) <= loadKernelChannel_CP_676_elements(11);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	43 
    -- CP-element group 18: 	44 
    -- CP-element group 18: 	65 
    -- CP-element group 18: 	64 
    -- CP-element group 18: 	86 
    -- CP-element group 18: 	24 
    -- CP-element group 18: 	25 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/$entry
      -- CP-element group 18: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/loop_body_start
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group loadKernelChannel_CP_676_elements(18) is bound as output of CP function.
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	86 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	29 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/condition_evaluated
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:do_while_stmt_349_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(19), ack => do_while_stmt_349_branch_req_0); -- 
    loadKernelChannel_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(86) & loadKernelChannel_CP_676_elements(23) & loadKernelChannel_CP_676_elements(29);
      gj_loadKernelChannel_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	43 
    -- CP-element group 20: 	24 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	26 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_sample_start__ps
      -- CP-element group 20: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/aggregated_phi_sample_req
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(20) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(43) & loadKernelChannel_CP_676_elements(24) & loadKernelChannel_CP_676_elements(23);
      gj_loadKernelChannel_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	45 
    -- CP-element group 21: 	27 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	75 
    -- CP-element group 21: 	79 
    -- CP-element group 21: 	83 
    -- CP-element group 21: 	87 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	43 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/aggregated_phi_sample_ack
      -- CP-element group 21: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_sample_completed_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(45) & loadKernelChannel_CP_676_elements(27);
      gj_loadKernelChannel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	44 
    -- CP-element group 22: 	25 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	28 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/aggregated_phi_update_req
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(22) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(44) & loadKernelChannel_CP_676_elements(25);
      gj_loadKernelChannel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	46 
    -- CP-element group 23: 	29 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(23) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(29);
      gj_loadKernelChannel_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_sample_start_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(21);
      gj_loadKernelChannel_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	72 
    -- CP-element group 25: 	80 
    -- CP-element group 25: 	66 
    -- CP-element group 25: 	61 
    -- CP-element group 25: 	29 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_update_start_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(72) & loadKernelChannel_CP_676_elements(80) & loadKernelChannel_CP_676_elements(66) & loadKernelChannel_CP_676_elements(61) & loadKernelChannel_CP_676_elements(29);
      gj_loadKernelChannel_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	20 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_sample_start__ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(26) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_CP_676_elements(26) <= loadKernelChannel_CP_676_elements(20);
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	21 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_sample_completed__ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(27) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group loadKernelChannel_CP_676_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	22 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_update_start__ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(28) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_CP_676_elements(28) <= loadKernelChannel_CP_676_elements(22);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	70 
    -- CP-element group 29: 	78 
    -- CP-element group 29: 	66 
    -- CP-element group 29: 	60 
    -- CP-element group 29: 	23 
    -- CP-element group 29: 	19 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (15) 
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_index_resize_1/index_resize_ack
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_index_resized_1
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_index_scale_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_index_scale_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_index_computed_1
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_index_scale_1/scale_rename_req
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_index_resize_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_index_resize_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_index_scale_1/scale_rename_ack
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_final_index_sum_regn_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_index_resize_1/index_resize_req
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_final_index_sum_regn_Sample/req
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_index_scaled_1
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_update_completed__ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:array_obj_ref_396_index_offset_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(29), ack => array_obj_ref_396_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	16 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_loopback_trigger
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(30) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_CP_676_elements(30) <= loadKernelChannel_CP_676_elements(16);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_loopback_sample_req
      -- CP-element group 31: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_loopback_sample_req_ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:phi_stmt_351_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_351_loopback_sample_req_828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_351_loopback_sample_req_828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(31), ack => phi_stmt_351_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(31) is bound as output of CP function.
    -- CP-element group 32:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	17 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_entry_trigger
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(32) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_CP_676_elements(32) <= loadKernelChannel_CP_676_elements(17);
    -- CP-element group 33:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_entry_sample_req
      -- CP-element group 33: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_entry_sample_req_ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:phi_stmt_351_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_351_entry_sample_req_831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_351_entry_sample_req_831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(33), ack => phi_stmt_351_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_phi_mux_ack
      -- CP-element group 34: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_351_phi_mux_ack_ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:phi_stmt_351_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_351_phi_mux_ack_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_351_ack_0, ack => loadKernelChannel_CP_676_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_sample_start__ps
      -- CP-element group 35: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_Sample/req
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:nmycount_373_353_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(35), ack => nmycount_373_353_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_update_start__ps
      -- CP-element group 36: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_update_start_
      -- CP-element group 36: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_Update/req
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:nmycount_373_353_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(36), ack => nmycount_373_353_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_sample_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_Sample/ack
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:nmycount_373_353_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_373_353_buf_ack_0, ack => loadKernelChannel_CP_676_elements(37)); -- 
    -- CP-element group 38:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_update_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nmycount_353_Update/ack
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:nmycount_373_353_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_373_353_buf_ack_1, ack => loadKernelChannel_CP_676_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_Sample/req
      -- CP-element group 39: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_sample_start__ps
      -- CP-element group 39: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_sample_start_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:start_add_354_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(39), ack => start_add_354_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_Update/req
      -- CP-element group 40: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_update_start_
      -- CP-element group 40: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_update_start__ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:start_add_354_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(40), ack => start_add_354_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(40) is bound as output of CP function.
    -- CP-element group 41:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (4) 
      -- CP-element group 41: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_Sample/ack
      -- CP-element group 41: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_sample_completed__ps
      -- CP-element group 41: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_sample_completed_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:start_add_354_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_354_buf_ack_0, ack => loadKernelChannel_CP_676_elements(41)); -- 
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (4) 
      -- CP-element group 42: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_start_add_354_update_completed__ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:start_add_354_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_354_buf_ack_1, ack => loadKernelChannel_CP_676_elements(42)); -- 
    -- CP-element group 43:  join  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	18 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	77 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	85 
    -- CP-element group 43: 	21 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	20 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_sample_start_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(43) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(77) & loadKernelChannel_CP_676_elements(81) & loadKernelChannel_CP_676_elements(85) & loadKernelChannel_CP_676_elements(21);
      gj_loadKernelChannel_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	18 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: 	61 
    -- CP-element group 44: 	84 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	22 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_update_start_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(44) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(61) & loadKernelChannel_CP_676_elements(84);
      gj_loadKernelChannel_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	21 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_sample_completed__ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(45) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group loadKernelChannel_CP_676_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	60 
    -- CP-element group 46: 	82 
    -- CP-element group 46: 	23 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_update_completed__ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(46) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group loadKernelChannel_CP_676_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_loopback_trigger
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(47) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_CP_676_elements(47) <= loadKernelChannel_CP_676_elements(16);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_loopback_sample_req_ps
      -- CP-element group 48: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_loopback_sample_req
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:phi_stmt_355_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_355_loopback_sample_req_882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_355_loopback_sample_req_882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(48), ack => phi_stmt_355_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_entry_trigger
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(49) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_CP_676_elements(49) <= loadKernelChannel_CP_676_elements(17);
    -- CP-element group 50:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_entry_sample_req
      -- CP-element group 50: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_entry_sample_req_ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:phi_stmt_355_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_355_entry_sample_req_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_355_entry_sample_req_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(50), ack => phi_stmt_355_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_phi_mux_ack
      -- CP-element group 51: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/phi_stmt_355_phi_mux_ack_ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:phi_stmt_355_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_355_phi_mux_ack_888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_355_ack_0, ack => loadKernelChannel_CP_676_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_Sample/$entry
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:nfetch_val_418_357_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(52), ack => nfetch_val_418_357_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_Update/req
      -- CP-element group 53: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_update_start_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:nfetch_val_418_357_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(53), ack => nfetch_val_418_357_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_sample_completed_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:nfetch_val_418_357_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_418_357_buf_ack_0, ack => loadKernelChannel_CP_676_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_nfetch_val_357_update_completed_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:nfetch_val_418_357_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_418_357_buf_ack_1, ack => loadKernelChannel_CP_676_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_sample_start__ps
      -- CP-element group 56: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_Sample/$entry
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:my_fetch_338_358_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(56), ack => my_fetch_338_358_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_update_start_
      -- CP-element group 57: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_Update/req
      -- CP-element group 57: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_update_start__ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:my_fetch_338_358_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(57), ack => my_fetch_338_358_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_sample_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_Sample/ack
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:my_fetch_338_358_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_338_358_buf_ack_0, ack => loadKernelChannel_CP_676_elements(58)); -- 
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_Update/ack
      -- CP-element group 59: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/R_my_fetch_358_update_completed__ps
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:my_fetch_338_358_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_338_358_buf_ack_1, ack => loadKernelChannel_CP_676_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	46 
    -- CP-element group 60: 	29 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/WPIPE_kernel_pipe1_380_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/WPIPE_kernel_pipe1_380_Sample/req
      -- CP-element group 60: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/WPIPE_kernel_pipe1_380_Sample/$entry
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:WPIPE_kernel_pipe1_380_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(60), ack => WPIPE_kernel_pipe1_380_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(29) & loadKernelChannel_CP_676_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	44 
    -- CP-element group 61: 	25 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/WPIPE_kernel_pipe1_380_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/WPIPE_kernel_pipe1_380_update_start_
      -- CP-element group 61: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/WPIPE_kernel_pipe1_380_Update/req
      -- CP-element group 61: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/WPIPE_kernel_pipe1_380_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/WPIPE_kernel_pipe1_380_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/WPIPE_kernel_pipe1_380_Sample/$exit
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:WPIPE_kernel_pipe1_380_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:WPIPE_kernel_pipe1_380_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_380_inst_ack_0, ack => loadKernelChannel_CP_676_elements(61)); -- 
    req_939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(61), ack => WPIPE_kernel_pipe1_380_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	87 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/WPIPE_kernel_pipe1_380_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/WPIPE_kernel_pipe1_380_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/WPIPE_kernel_pipe1_380_Update/$exit
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:WPIPE_kernel_pipe1_380_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_380_inst_ack_1, ack => loadKernelChannel_CP_676_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	67 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	68 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	68 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/addr_of_397_request/$entry
      -- CP-element group 63: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/addr_of_397_request/req
      -- CP-element group 63: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/addr_of_397_sample_start_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:addr_of_397_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(63), ack => addr_of_397_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(67) & loadKernelChannel_CP_676_elements(68);
      gj_loadKernelChannel_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	18 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	76 
    -- CP-element group 64: 	69 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/addr_of_397_complete/$entry
      -- CP-element group 64: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/addr_of_397_complete/req
      -- CP-element group 64: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/addr_of_397_update_start_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:addr_of_397_final_reg_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(64), ack => addr_of_397_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(76) & loadKernelChannel_CP_676_elements(69);
      gj_loadKernelChannel_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	68 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_final_index_sum_regn_Update/req
      -- CP-element group 65: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_final_index_sum_regn_update_start
      -- CP-element group 65: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_final_index_sum_regn_Update/$entry
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:array_obj_ref_396_index_offset_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(65), ack => array_obj_ref_396_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(67) & loadKernelChannel_CP_676_elements(68);
      gj_loadKernelChannel_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	29 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	87 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	25 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_final_index_sum_regn_sample_complete
      -- CP-element group 66: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_final_index_sum_regn_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:array_obj_ref_396_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_396_index_offset_ack_0, ack => loadKernelChannel_CP_676_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	63 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (8) 
      -- CP-element group 67: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_final_index_sum_regn_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_final_index_sum_regn_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_offset_calculated
      -- CP-element group 67: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_base_plus_offset/$entry
      -- CP-element group 67: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_base_plus_offset/$exit
      -- CP-element group 67: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_base_plus_offset/sum_rename_req
      -- CP-element group 67: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_base_plus_offset/sum_rename_ack
      -- CP-element group 67: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/array_obj_ref_396_root_address_calculated
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:array_obj_ref_396_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_396_index_offset_ack_1, ack => loadKernelChannel_CP_676_elements(67)); -- 
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	63 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	63 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/addr_of_397_request/$exit
      -- CP-element group 68: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/addr_of_397_request/ack
      -- CP-element group 68: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/addr_of_397_sample_completed_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:addr_of_397_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_397_final_reg_ack_0, ack => loadKernelChannel_CP_676_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	64 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	64 
    -- CP-element group 69:  members (19) 
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_base_addr_resize/base_resize_req
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_root_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_word_addrgen/root_register_ack
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_base_plus_offset/sum_rename_req
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_word_addrgen/$entry
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_base_plus_offset/$exit
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_base_plus_offset/sum_rename_ack
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/addr_of_397_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_word_addrgen/$exit
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_base_addr_resize/$exit
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/addr_of_397_complete/$exit
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/addr_of_397_complete/ack
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_base_addr_resize/base_resize_ack
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_base_address_resized
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_word_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_base_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_base_addr_resize/$entry
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_base_plus_offset/$entry
      -- CP-element group 69: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_word_addrgen/root_register_req
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:addr_of_397_final_reg_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_397_final_reg_ack_1, ack => loadKernelChannel_CP_676_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	29 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_401_Sample/req
      -- CP-element group 70: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_401_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_401_Sample/$entry
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(70) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:W_fn_387_delayed_7_0_399_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(70), ack => W_fn_387_delayed_7_0_399_inst_req_0); -- 
    loadKernelChannel_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(29) & loadKernelChannel_CP_676_elements(72);
      gj_loadKernelChannel_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	76 
    -- CP-element group 71: 	73 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_401_update_start_
      -- CP-element group 71: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_401_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_401_Update/req
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(71) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:W_fn_387_delayed_7_0_399_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(71), ack => W_fn_387_delayed_7_0_399_inst_req_1); -- 
    loadKernelChannel_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(76) & loadKernelChannel_CP_676_elements(73);
      gj_loadKernelChannel_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	25 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_401_Sample/ack
      -- CP-element group 72: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_401_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_401_Sample/$exit
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(72) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:W_fn_387_delayed_7_0_399_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_387_delayed_7_0_399_inst_ack_0, ack => loadKernelChannel_CP_676_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_401_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_401_Update/ack
      -- CP-element group 73: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_401_Update/$exit
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:W_fn_387_delayed_7_0_399_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_387_delayed_7_0_399_inst_ack_1, ack => loadKernelChannel_CP_676_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: 	69 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Sample/word_access_start/word_0/rr
      -- CP-element group 74: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Sample/word_access_start/word_0/$entry
      -- CP-element group 74: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Sample/word_access_start/$entry
      -- CP-element group 74: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Sample/$entry
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:ptr_deref_405_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(74), ack => ptr_deref_405_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(73) & loadKernelChannel_CP_676_elements(69) & loadKernelChannel_CP_676_elements(76);
      gj_loadKernelChannel_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	21 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_update_start_
      -- CP-element group 75: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Update/word_access_complete/word_0/cr
      -- CP-element group 75: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Update/word_access_complete/word_0/$entry
      -- CP-element group 75: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Update/word_access_complete/$entry
      -- CP-element group 75: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Update/$entry
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:ptr_deref_405_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(75), ack => ptr_deref_405_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(77);
      gj_loadKernelChannel_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	71 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	64 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Sample/word_access_start/word_0/ra
      -- CP-element group 76: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Sample/word_access_start/word_0/$exit
      -- CP-element group 76: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Sample/word_access_start/$exit
      -- CP-element group 76: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Sample/$exit
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:ptr_deref_405_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_405_load_0_ack_0, ack => loadKernelChannel_CP_676_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	87 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	43 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Update/ptr_deref_405_Merge/$entry
      -- CP-element group 77: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Update/word_access_complete/word_0/ca
      -- CP-element group 77: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Update/ptr_deref_405_Merge/merge_req
      -- CP-element group 77: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Update/ptr_deref_405_Merge/merge_ack
      -- CP-element group 77: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Update/ptr_deref_405_Merge/$exit
      -- CP-element group 77: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Update/word_access_complete/word_0/$exit
      -- CP-element group 77: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Update/word_access_complete/$exit
      -- CP-element group 77: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/ptr_deref_405_Update/$exit
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:ptr_deref_405_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_405_load_0_ack_1, ack => loadKernelChannel_CP_676_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	29 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_409_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_409_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_409_Sample/req
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(78) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:W_fn_393_delayed_13_0_407_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(78), ack => W_fn_393_delayed_13_0_407_inst_req_0); -- 
    loadKernelChannel_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(29) & loadKernelChannel_CP_676_elements(80);
      gj_loadKernelChannel_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	21 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	81 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_409_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_409_Update/req
      -- CP-element group 79: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_409_update_start_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:W_fn_393_delayed_13_0_407_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(79), ack => W_fn_393_delayed_13_0_407_inst_req_1); -- 
    loadKernelChannel_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(81);
      gj_loadKernelChannel_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	25 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_409_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_409_Sample/ack
      -- CP-element group 80: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_409_Sample/$exit
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:W_fn_393_delayed_13_0_407_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_393_delayed_13_0_407_inst_ack_0, ack => loadKernelChannel_CP_676_elements(80)); -- 
    -- CP-element group 81:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	87 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	43 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_409_Update/ack
      -- CP-element group 81: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_409_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_409_update_completed_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(81) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:W_fn_393_delayed_13_0_407_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_393_delayed_13_0_407_inst_ack_1, ack => loadKernelChannel_CP_676_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	46 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_412_Sample/req
      -- CP-element group 82: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_412_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_412_sample_start_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:W_fetch_val_395_delayed_13_0_410_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(82), ack => W_fetch_val_395_delayed_13_0_410_inst_req_0); -- 
    loadKernelChannel_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(84);
      gj_loadKernelChannel_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	21 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_412_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_412_Update/req
      -- CP-element group 83: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_412_update_start_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(83) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:W_fetch_val_395_delayed_13_0_410_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(83), ack => W_fetch_val_395_delayed_13_0_410_inst_req_1); -- 
    loadKernelChannel_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(85);
      gj_loadKernelChannel_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	44 
    -- CP-element group 84: 	82 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_412_Sample/ack
      -- CP-element group 84: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_412_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_412_sample_completed_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(84) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:W_fetch_val_395_delayed_13_0_410_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_395_delayed_13_0_410_inst_ack_0, ack => loadKernelChannel_CP_676_elements(84)); -- 
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	43 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_412_Update/ack
      -- CP-element group 85: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_412_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/assign_stmt_412_update_completed_
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(85) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:W_fetch_val_395_delayed_13_0_410_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_395_delayed_13_0_410_inst_ack_1, ack => loadKernelChannel_CP_676_elements(85)); -- 
    -- CP-element group 86:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	18 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	19 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(86) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group loadKernelChannel_CP_676_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_676_elements(18), ack => loadKernelChannel_CP_676_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	77 
    -- CP-element group 87: 	66 
    -- CP-element group 87: 	62 
    -- CP-element group 87: 	81 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	21 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	15 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_348/do_while_stmt_349/do_while_stmt_349_loop_body/$exit
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(87) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(77) & loadKernelChannel_CP_676_elements(66) & loadKernelChannel_CP_676_elements(62) & loadKernelChannel_CP_676_elements(81) & loadKernelChannel_CP_676_elements(85) & loadKernelChannel_CP_676_elements(21);
      gj_loadKernelChannel_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	14 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_348/do_while_stmt_349/loop_exit/$exit
      -- CP-element group 88: 	 branch_block_stmt_348/do_while_stmt_349/loop_exit/ack
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:do_while_stmt_349_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_349_branch_ack_0, ack => loadKernelChannel_CP_676_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	14 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_348/do_while_stmt_349/loop_taken/ack
      -- CP-element group 89: 	 branch_block_stmt_348/do_while_stmt_349/loop_taken/$exit
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:do_while_stmt_349_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_349_branch_ack_1, ack => loadKernelChannel_CP_676_elements(89)); -- 
    -- CP-element group 90:  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	12 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	10 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_348/do_while_stmt_349/$exit
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(90) fired."); 
        -- 
      end if; --
    end process; 
    loadKernelChannel_CP_676_elements(90) <= loadKernelChannel_CP_676_elements(12);
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	10 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 assign_stmt_432/type_cast_431_sample_completed_
      -- CP-element group 91: 	 assign_stmt_432/type_cast_431_Sample/$exit
      -- CP-element group 91: 	 assign_stmt_432/type_cast_431_Sample/ra
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(91) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:type_cast_431_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_431_inst_ack_0, ack => loadKernelChannel_CP_676_elements(91)); -- 
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	10 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 assign_stmt_432/WPIPE_size_pipe_427_Sample/req
      -- CP-element group 92: 	 assign_stmt_432/type_cast_431_update_completed_
      -- CP-element group 92: 	 assign_stmt_432/WPIPE_size_pipe_427_sample_start_
      -- CP-element group 92: 	 assign_stmt_432/type_cast_431_Update/ca
      -- CP-element group 92: 	 assign_stmt_432/type_cast_431_Update/$exit
      -- CP-element group 92: 	 assign_stmt_432/WPIPE_size_pipe_427_Sample/$entry
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(92) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:type_cast_431_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:WPIPE_size_pipe_427_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_431_inst_ack_1, ack => loadKernelChannel_CP_676_elements(92)); -- 
    req_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(92), ack => WPIPE_size_pipe_427_inst_req_0); -- 
    -- CP-element group 93:  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 assign_stmt_432/WPIPE_size_pipe_427_update_start_
      -- CP-element group 93: 	 assign_stmt_432/WPIPE_size_pipe_427_Update/req
      -- CP-element group 93: 	 assign_stmt_432/WPIPE_size_pipe_427_Sample/$exit
      -- CP-element group 93: 	 assign_stmt_432/WPIPE_size_pipe_427_sample_completed_
      -- CP-element group 93: 	 assign_stmt_432/WPIPE_size_pipe_427_Update/$entry
      -- CP-element group 93: 	 assign_stmt_432/WPIPE_size_pipe_427_Sample/ack
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:WPIPE_size_pipe_427_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:WPIPE_size_pipe_427_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_427_inst_ack_0, ack => loadKernelChannel_CP_676_elements(93)); -- 
    req_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(93), ack => WPIPE_size_pipe_427_inst_req_1); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 assign_stmt_432/WPIPE_size_pipe_427_update_completed_
      -- CP-element group 94: 	 assign_stmt_432/WPIPE_size_pipe_427_Update/ack
      -- CP-element group 94: 	 assign_stmt_432/WPIPE_size_pipe_427_Update/$exit
      -- CP-element group 94: 	 $exit
      -- CP-element group 94: 	 assign_stmt_432/$exit
      -- 
    -- logger for CP element group loadKernelChannel_CP_676_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadKernelChannel_CP_676_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:loadKernelChannel_CP_676_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadKernelChannel:CP:WPIPE_size_pipe_427_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_427_inst_ack_1, ack => loadKernelChannel_CP_676_elements(94)); -- 
    loadKernelChannel_do_while_stmt_349_terminator_1088: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_349_terminator_1088", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_676_elements(15),loop_continue => loadKernelChannel_CP_676_elements(89),loop_terminate => loadKernelChannel_CP_676_elements(88),loop_back => loadKernelChannel_CP_676_elements(13),loop_exit => loadKernelChannel_CP_676_elements(12),clk => clk, reset => reset); -- 
    phi_stmt_351_phi_seq_872_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_676_elements(30);
      loadKernelChannel_CP_676_elements(35)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_676_elements(37);
      loadKernelChannel_CP_676_elements(36)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_676_elements(38);
      loadKernelChannel_CP_676_elements(31) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_676_elements(32);
      loadKernelChannel_CP_676_elements(39)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_676_elements(41);
      loadKernelChannel_CP_676_elements(40)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_676_elements(42);
      loadKernelChannel_CP_676_elements(33) <= phi_mux_reqs(1);
      phi_stmt_351_phi_seq_872 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_351_phi_seq_872") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_676_elements(26), 
          phi_sample_ack => loadKernelChannel_CP_676_elements(27), 
          phi_update_req => loadKernelChannel_CP_676_elements(28), 
          phi_update_ack => loadKernelChannel_CP_676_elements(29), 
          phi_mux_ack => loadKernelChannel_CP_676_elements(34), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_355_phi_seq_926_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_676_elements(47);
      loadKernelChannel_CP_676_elements(52)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_676_elements(54);
      loadKernelChannel_CP_676_elements(53)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_676_elements(55);
      loadKernelChannel_CP_676_elements(48) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_676_elements(49);
      loadKernelChannel_CP_676_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_676_elements(58);
      loadKernelChannel_CP_676_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_676_elements(59);
      loadKernelChannel_CP_676_elements(50) <= phi_mux_reqs(1);
      phi_stmt_355_phi_seq_926 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_355_phi_seq_926") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_676_elements(20), 
          phi_sample_ack => loadKernelChannel_CP_676_elements(45), 
          phi_update_req => loadKernelChannel_CP_676_elements(22), 
          phi_update_ack => loadKernelChannel_CP_676_elements(46), 
          phi_mux_ack => loadKernelChannel_CP_676_elements(51), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_814_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_676_elements(16);
        preds(1)  <= loadKernelChannel_CP_676_elements(17);
        entry_tmerge_814 : transition_merge -- 
          generic map(name => " entry_tmerge_814")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_676_elements(18));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u64_u64_364_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_386_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_377_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_395_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_395_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_395_wire : std_logic_vector(63 downto 0);
    signal R_sh_start_331_resized : std_logic_vector(13 downto 0);
    signal R_sh_start_331_scaled : std_logic_vector(13 downto 0);
    signal SUB_u64_u64_365_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_423_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_430_wire : std_logic_vector(63 downto 0);
    signal ULT_u64_u1_424_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_332_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_332_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_332_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_332_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_332_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_332_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_396_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_396_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_396_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_396_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_396_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_396_root_address : std_logic_vector(13 downto 0);
    signal fetch_addr_334 : std_logic_vector(31 downto 0);
    signal fetch_addr_398 : std_logic_vector(31 downto 0);
    signal fetch_val_355 : std_logic_vector(63 downto 0);
    signal fetch_val_395_delayed_13_0_412 : std_logic_vector(63 downto 0);
    signal first_fill_343 : std_logic_vector(0 downto 0);
    signal fn_387_delayed_7_0_401 : std_logic_vector(0 downto 0);
    signal fn_389 : std_logic_vector(0 downto 0);
    signal fn_393_delayed_13_0_409 : std_logic_vector(0 downto 0);
    signal fv_406 : std_logic_vector(63 downto 0);
    signal konst_325_wire_constant : std_logic_vector(63 downto 0);
    signal konst_341_wire_constant : std_logic_vector(63 downto 0);
    signal konst_361_wire_constant : std_logic_vector(63 downto 0);
    signal konst_363_wire_constant : std_logic_vector(63 downto 0);
    signal konst_366_wire_constant : std_logic_vector(63 downto 0);
    signal konst_371_wire_constant : std_logic_vector(63 downto 0);
    signal konst_385_wire_constant : std_logic_vector(63 downto 0);
    signal konst_387_wire_constant : std_logic_vector(63 downto 0);
    signal konst_394_wire_constant : std_logic_vector(63 downto 0);
    signal konst_422_wire_constant : std_logic_vector(63 downto 0);
    signal my_fetch_338 : std_logic_vector(63 downto 0);
    signal my_fetch_338_358_buffered : std_logic_vector(63 downto 0);
    signal my_num1_368 : std_logic_vector(63 downto 0);
    signal mycount_351 : std_logic_vector(63 downto 0);
    signal nfetch_val_418 : std_logic_vector(63 downto 0);
    signal nfetch_val_418_357_buffered : std_logic_vector(63 downto 0);
    signal nmycount_373 : std_logic_vector(63 downto 0);
    signal nmycount_373_353_buffered : std_logic_vector(63 downto 0);
    signal ptr_deref_337_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_337_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_337_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_337_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_337_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_405_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_405_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_405_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_405_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_405_word_offset_0 : std_logic_vector(13 downto 0);
    signal sh_start_327 : std_logic_vector(63 downto 0);
    signal start_add_354_buffered : std_logic_vector(63 downto 0);
    signal start_next_347 : std_logic_vector(0 downto 0);
    signal type_cast_431_wire : std_logic_vector(31 downto 0);
    signal var_val_379 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_332_constant_part_of_offset <= "00000000000000";
    array_obj_ref_332_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_332_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_332_resized_base_address <= "00000000000000";
    array_obj_ref_396_constant_part_of_offset <= "00000000000000";
    array_obj_ref_396_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_396_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_396_resized_base_address <= "00000000000000";
    konst_325_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_341_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_361_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_363_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_366_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_371_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_385_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_387_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_394_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_422_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    ptr_deref_337_word_offset_0 <= "00000000000000";
    ptr_deref_405_word_offset_0 <= "00000000000000";
    -- logger for phi phi_stmt_351
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_351_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:loadKernelChannel:DP:phi_stmt_351:input-0 nmycount_373_353_buffered= " & Convert_SLV_To_Hex_String(nmycount_373_353_buffered));
          --
        end if;
        if phi_stmt_351_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:loadKernelChannel:DP:phi_stmt_351:input-1 start_add_354_buffered= " & Convert_SLV_To_Hex_String(start_add_354_buffered));
          --
        end if;
        if phi_stmt_351_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:loadKernelChannel:DP:phi_stmt_351:sample-completed");
          --
        end if;
        if phi_stmt_351_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:loadKernelChannel:DP:phi_stmt_351:output mycount_351= " & Convert_SLV_To_Hex_String(mycount_351));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_351: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_373_353_buffered & start_add_354_buffered;
      req <= phi_stmt_351_req_0 & phi_stmt_351_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_351",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_351_ack_0,
          idata => idata,
          odata => mycount_351,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_351
    -- logger for phi phi_stmt_355
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_355_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:loadKernelChannel:DP:phi_stmt_355:input-0 nfetch_val_418_357_buffered= " & Convert_SLV_To_Hex_String(nfetch_val_418_357_buffered));
          --
        end if;
        if phi_stmt_355_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:loadKernelChannel:DP:phi_stmt_355:input-1 my_fetch_338_358_buffered= " & Convert_SLV_To_Hex_String(my_fetch_338_358_buffered));
          --
        end if;
        if phi_stmt_355_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:loadKernelChannel:DP:phi_stmt_355:sample-completed");
          --
        end if;
        if phi_stmt_355_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:loadKernelChannel:DP:phi_stmt_355:output fetch_val_355= " & Convert_SLV_To_Hex_String(fetch_val_355));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_355: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nfetch_val_418_357_buffered & my_fetch_338_358_buffered;
      req <= phi_stmt_355_req_0 & phi_stmt_355_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_355",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_355_ack_0,
          idata => idata,
          odata => fetch_val_355,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_355
    -- logger for split-operator MUX_417_inst flow-through 
    process(nfetch_val_418) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:MUX_417_inst:flowthrough inputs: " & " fn_393_delayed_13_0_409 = "& Convert_SLV_To_Hex_String(fn_393_delayed_13_0_409) & " fv_406 = "& Convert_SLV_To_Hex_String(fv_406) & " fetch_val_395_delayed_13_0_412 = "& Convert_SLV_To_Hex_String(fetch_val_395_delayed_13_0_412) & " outputs:" & " nfetch_val_418= "  & Convert_SLV_To_Hex_String(nfetch_val_418));
      --
    end process; 
    -- flow-through select operator MUX_417_inst
    nfetch_val_418 <= fv_406 when (fn_393_delayed_13_0_409(0) /=  '0') else fetch_val_395_delayed_13_0_412;
    -- logger for split-operator W_fetch_val_395_delayed_13_0_410_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_fetch_val_395_delayed_13_0_410_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:W_fetch_val_395_delayed_13_0_410_inst:started:   inputs: " & " fetch_val_355 = "& Convert_SLV_To_Hex_String(fetch_val_355));
          --
        end if; 
        if W_fetch_val_395_delayed_13_0_410_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:W_fetch_val_395_delayed_13_0_410_inst:finished:  outputs: " & " fetch_val_395_delayed_13_0_412= "  & Convert_SLV_To_Hex_String(fetch_val_395_delayed_13_0_412));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_fetch_val_395_delayed_13_0_410_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val_395_delayed_13_0_410_inst_req_0;
      W_fetch_val_395_delayed_13_0_410_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val_395_delayed_13_0_410_inst_req_1;
      W_fetch_val_395_delayed_13_0_410_inst_ack_1<= rack(0);
      W_fetch_val_395_delayed_13_0_410_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val_395_delayed_13_0_410_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val_355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val_395_delayed_13_0_412,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_fn_387_delayed_7_0_399_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_fn_387_delayed_7_0_399_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:W_fn_387_delayed_7_0_399_inst:started:   inputs: " & " fn_389 = "& Convert_SLV_To_Hex_String(fn_389));
          --
        end if; 
        if W_fn_387_delayed_7_0_399_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:W_fn_387_delayed_7_0_399_inst:finished:  outputs: " & " fn_387_delayed_7_0_401= "  & Convert_SLV_To_Hex_String(fn_387_delayed_7_0_401));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_fn_387_delayed_7_0_399_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_387_delayed_7_0_399_inst_req_0;
      W_fn_387_delayed_7_0_399_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_387_delayed_7_0_399_inst_req_1;
      W_fn_387_delayed_7_0_399_inst_ack_1<= rack(0);
      W_fn_387_delayed_7_0_399_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_387_delayed_7_0_399_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_389,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_387_delayed_7_0_401,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_fn_393_delayed_13_0_407_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_fn_393_delayed_13_0_407_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:W_fn_393_delayed_13_0_407_inst:started:   inputs: " & " fn_389 = "& Convert_SLV_To_Hex_String(fn_389));
          --
        end if; 
        if W_fn_393_delayed_13_0_407_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:W_fn_393_delayed_13_0_407_inst:finished:  outputs: " & " fn_393_delayed_13_0_409= "  & Convert_SLV_To_Hex_String(fn_393_delayed_13_0_409));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_fn_393_delayed_13_0_407_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_393_delayed_13_0_407_inst_req_0;
      W_fn_393_delayed_13_0_407_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_393_delayed_13_0_407_inst_req_1;
      W_fn_393_delayed_13_0_407_inst_ack_1<= rack(0);
      W_fn_393_delayed_13_0_407_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_393_delayed_13_0_407_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_389,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_393_delayed_13_0_409,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_333_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_333_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:addr_of_333_final_reg:started:   inputs: " & " array_obj_ref_332_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_332_root_address));
          --
        end if; 
        if addr_of_333_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:addr_of_333_final_reg:finished:  outputs: " & " fetch_addr_334= "  & Convert_SLV_To_Hex_String(fetch_addr_334));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_333_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_333_final_reg_req_0;
      addr_of_333_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_333_final_reg_req_1;
      addr_of_333_final_reg_ack_1<= rack(0);
      addr_of_333_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_333_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_332_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_334,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_397_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_397_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:addr_of_397_final_reg:started:   inputs: " & " array_obj_ref_396_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_396_root_address));
          --
        end if; 
        if addr_of_397_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:addr_of_397_final_reg:finished:  outputs: " & " fetch_addr_398= "  & Convert_SLV_To_Hex_String(fetch_addr_398));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_397_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_397_final_reg_req_0;
      addr_of_397_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_397_final_reg_req_1;
      addr_of_397_final_reg_ack_1<= rack(0);
      addr_of_397_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_397_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_396_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_398,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator my_fetch_338_358_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if my_fetch_338_358_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:my_fetch_338_358_buf:started:   inputs: " & " my_fetch_338 = "& Convert_SLV_To_Hex_String(my_fetch_338));
          --
        end if; 
        if my_fetch_338_358_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:my_fetch_338_358_buf:finished:  outputs: " & " my_fetch_338_358_buffered= "  & Convert_SLV_To_Hex_String(my_fetch_338_358_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    my_fetch_338_358_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch_338_358_buf_req_0;
      my_fetch_338_358_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch_338_358_buf_req_1;
      my_fetch_338_358_buf_ack_1<= rack(0);
      my_fetch_338_358_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch_338_358_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch_338,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch_338_358_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator nfetch_val_418_357_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if nfetch_val_418_357_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:nfetch_val_418_357_buf:started:   inputs: " & " nfetch_val_418 = "& Convert_SLV_To_Hex_String(nfetch_val_418));
          --
        end if; 
        if nfetch_val_418_357_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:nfetch_val_418_357_buf:finished:  outputs: " & " nfetch_val_418_357_buffered= "  & Convert_SLV_To_Hex_String(nfetch_val_418_357_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    nfetch_val_418_357_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nfetch_val_418_357_buf_req_0;
      nfetch_val_418_357_buf_ack_0<= wack(0);
      rreq(0) <= nfetch_val_418_357_buf_req_1;
      nfetch_val_418_357_buf_ack_1<= rack(0);
      nfetch_val_418_357_buf : InterlockBuffer generic map ( -- 
        name => "nfetch_val_418_357_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nfetch_val_418,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nfetch_val_418_357_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator nmycount_373_353_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if nmycount_373_353_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:nmycount_373_353_buf:started:   inputs: " & " nmycount_373 = "& Convert_SLV_To_Hex_String(nmycount_373));
          --
        end if; 
        if nmycount_373_353_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:nmycount_373_353_buf:finished:  outputs: " & " nmycount_373_353_buffered= "  & Convert_SLV_To_Hex_String(nmycount_373_353_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    nmycount_373_353_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_373_353_buf_req_0;
      nmycount_373_353_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_373_353_buf_req_1;
      nmycount_373_353_buf_ack_1<= rack(0);
      nmycount_373_353_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_373_353_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_373,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_373_353_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator start_add_354_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if start_add_354_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:start_add_354_buf:started:   inputs: " & " start_add_buffer = "& Convert_SLV_To_Hex_String(start_add_buffer));
          --
        end if; 
        if start_add_354_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:start_add_354_buf:finished:  outputs: " & " start_add_354_buffered= "  & Convert_SLV_To_Hex_String(start_add_354_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    start_add_354_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_354_buf_req_0;
      start_add_354_buf_ack_0<= wack(0);
      rreq(0) <= start_add_354_buf_req_1;
      start_add_354_buf_ack_1<= rack(0);
      start_add_354_buf : InterlockBuffer generic map ( -- 
        name => "start_add_354_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_354_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_378_inst flow-through 
    process(var_val_379) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:type_cast_378_inst:flowthrough inputs: " & " LSHR_u64_u64_377_wire = "& Convert_SLV_To_Hex_String(LSHR_u64_u64_377_wire) & " outputs:" & " var_val_379= "  & Convert_SLV_To_Hex_String(var_val_379));
      --
    end process; 
    -- interlock type_cast_378_inst
    process(LSHR_u64_u64_377_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_377_wire(15 downto 0);
      var_val_379 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_431_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_431_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:type_cast_431_inst:started:   inputs: " & " first_fill_343 (guard)= " & Convert_SLV_To_String(first_fill_343) & " SUB_u64_u64_430_wire = "& Convert_SLV_To_Hex_String(SUB_u64_u64_430_wire));
          --
        end if; 
        if type_cast_431_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:type_cast_431_inst:finished:  outputs: " & " type_cast_431_wire= "  & Convert_SLV_To_Hex_String(type_cast_431_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_431_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_431_inst_req_0;
      type_cast_431_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_431_inst_req_1;
      type_cast_431_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  first_fill_343(0);
      type_cast_431_inst_gI: SplitGuardInterface generic map(name => "type_cast_431_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_431_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_431_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => SUB_u64_u64_430_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_431_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_332_index_1_rename flow-through 
    process(R_sh_start_331_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:array_obj_ref_332_index_1_rename:flowthrough  inputs: " & " R_sh_start_331_resized = "& Convert_SLV_To_Hex_String(R_sh_start_331_resized) & "outputs: " & " R_sh_start_331_scaled= "  & Convert_SLV_To_Hex_String(R_sh_start_331_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_332_index_1_rename
    process(R_sh_start_331_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_sh_start_331_resized;
      ov(13 downto 0) := iv;
      R_sh_start_331_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_332_index_1_resize flow-through 
    process(R_sh_start_331_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:array_obj_ref_332_index_1_resize:flowthrough  inputs: " & " sh_start_327 = "& Convert_SLV_To_Hex_String(sh_start_327) & "outputs: " & " R_sh_start_331_resized= "  & Convert_SLV_To_Hex_String(R_sh_start_331_resized));
      --
    end process; 
    -- equivalence array_obj_ref_332_index_1_resize
    process(sh_start_327) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := sh_start_327;
      ov := iv(13 downto 0);
      R_sh_start_331_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_332_root_address_inst flow-through 
    process(array_obj_ref_332_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:array_obj_ref_332_root_address_inst:flowthrough  inputs: " & " array_obj_ref_332_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_332_final_offset) & "outputs: " & " array_obj_ref_332_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_332_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_332_root_address_inst
    process(array_obj_ref_332_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_332_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_332_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_396_index_1_rename flow-through 
    process(LSHR_u64_u64_395_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:array_obj_ref_396_index_1_rename:flowthrough  inputs: " & " LSHR_u64_u64_395_resized = "& Convert_SLV_To_Hex_String(LSHR_u64_u64_395_resized) & "outputs: " & " LSHR_u64_u64_395_scaled= "  & Convert_SLV_To_Hex_String(LSHR_u64_u64_395_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_396_index_1_rename
    process(LSHR_u64_u64_395_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_395_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_395_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_396_index_1_resize flow-through 
    process(LSHR_u64_u64_395_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:array_obj_ref_396_index_1_resize:flowthrough  inputs: " & " LSHR_u64_u64_395_wire = "& Convert_SLV_To_Hex_String(LSHR_u64_u64_395_wire) & "outputs: " & " LSHR_u64_u64_395_resized= "  & Convert_SLV_To_Hex_String(LSHR_u64_u64_395_resized));
      --
    end process; 
    -- equivalence array_obj_ref_396_index_1_resize
    process(LSHR_u64_u64_395_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_395_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_395_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_396_root_address_inst flow-through 
    process(array_obj_ref_396_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:array_obj_ref_396_root_address_inst:flowthrough  inputs: " & " array_obj_ref_396_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_396_final_offset) & "outputs: " & " array_obj_ref_396_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_396_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_396_root_address_inst
    process(array_obj_ref_396_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_396_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_396_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_337_addr_0 flow-through 
    process(ptr_deref_337_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ptr_deref_337_addr_0:flowthrough  inputs: " & " ptr_deref_337_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_337_root_address) & "outputs: " & " ptr_deref_337_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_337_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_337_addr_0
    process(ptr_deref_337_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_337_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_337_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_337_base_resize flow-through 
    process(ptr_deref_337_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ptr_deref_337_base_resize:flowthrough  inputs: " & " fetch_addr_334 = "& Convert_SLV_To_Hex_String(fetch_addr_334) & "outputs: " & " ptr_deref_337_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_337_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_337_base_resize
    process(fetch_addr_334) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_334;
      ov := iv(13 downto 0);
      ptr_deref_337_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_337_gather_scatter flow-through 
    process(my_fetch_338) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ptr_deref_337_gather_scatter:flowthrough  inputs: " & " ptr_deref_337_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_337_data_0) & "outputs: " & " my_fetch_338= "  & Convert_SLV_To_Hex_String(my_fetch_338));
      --
    end process; 
    -- equivalence ptr_deref_337_gather_scatter
    process(ptr_deref_337_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_337_data_0;
      ov(63 downto 0) := iv;
      my_fetch_338 <= ov(63 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_337_root_address_inst flow-through 
    process(ptr_deref_337_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ptr_deref_337_root_address_inst:flowthrough  inputs: " & " ptr_deref_337_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_337_resized_base_address) & "outputs: " & " ptr_deref_337_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_337_root_address));
      --
    end process; 
    -- equivalence ptr_deref_337_root_address_inst
    process(ptr_deref_337_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_337_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_337_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_405_addr_0 flow-through 
    process(ptr_deref_405_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ptr_deref_405_addr_0:flowthrough  inputs: " & " fn_387_delayed_7_0_401 (guard)= " & Convert_SLV_To_String(fn_387_delayed_7_0_401) & " ptr_deref_405_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_405_root_address) & "outputs: " & " ptr_deref_405_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_405_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_405_addr_0
    process(ptr_deref_405_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_405_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_405_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_405_base_resize flow-through 
    process(ptr_deref_405_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ptr_deref_405_base_resize:flowthrough  inputs: " & " fn_387_delayed_7_0_401 (guard)= " & Convert_SLV_To_String(fn_387_delayed_7_0_401) & " fetch_addr_398 = "& Convert_SLV_To_Hex_String(fetch_addr_398) & "outputs: " & " ptr_deref_405_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_405_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_405_base_resize
    process(fetch_addr_398) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_398;
      ov := iv(13 downto 0);
      ptr_deref_405_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_405_gather_scatter flow-through 
    process(fv_406) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ptr_deref_405_gather_scatter:flowthrough  inputs: " & " fn_387_delayed_7_0_401 (guard)= " & Convert_SLV_To_String(fn_387_delayed_7_0_401) & " ptr_deref_405_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_405_data_0) & "outputs: " & " fv_406= "  & Convert_SLV_To_Hex_String(fv_406));
      --
    end process; 
    -- equivalence ptr_deref_405_gather_scatter
    process(ptr_deref_405_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_405_data_0;
      ov(63 downto 0) := iv;
      fv_406 <= ov(63 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_405_root_address_inst flow-through 
    process(ptr_deref_405_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ptr_deref_405_root_address_inst:flowthrough  inputs: " & " fn_387_delayed_7_0_401 (guard)= " & Convert_SLV_To_String(fn_387_delayed_7_0_401) & " ptr_deref_405_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_405_resized_base_address) & "outputs: " & " ptr_deref_405_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_405_root_address));
      --
    end process; 
    -- equivalence ptr_deref_405_root_address_inst
    process(ptr_deref_405_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_405_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_405_root_address <= ov(13 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_349_branch_req_0," req0 do_while_stmt_349_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_349_branch_ack_0," ack0 do_while_stmt_349_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_349_branch_ack_1," ack1 do_while_stmt_349_branch");
    do_while_stmt_349_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u64_u1_424_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_349_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_349_branch_req_0,
          ack0 => do_while_stmt_349_branch_ack_0,
          ack1 => do_while_stmt_349_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u64_u64_372_inst flow-through 
    process(nmycount_373) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ADD_u64_u64_372_inst:flowthrough inputs: " & " mycount_351 = "& Convert_SLV_To_Hex_String(mycount_351) & " konst_371_wire_constant = "& Convert_SLV_To_Hex_String(konst_371_wire_constant) & " outputs:" & " nmycount_373= "  & Convert_SLV_To_Hex_String(nmycount_373));
      --
    end process; 
    -- binary operator ADD_u64_u64_372_inst
    process(mycount_351) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_351, konst_371_wire_constant, tmp_var);
      nmycount_373 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u64_u64_364_inst flow-through 
    process(AND_u64_u64_364_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:AND_u64_u64_364_inst:flowthrough inputs: " & " mycount_351 = "& Convert_SLV_To_Hex_String(mycount_351) & " konst_363_wire_constant = "& Convert_SLV_To_Hex_String(konst_363_wire_constant) & " outputs:" & " AND_u64_u64_364_wire= "  & Convert_SLV_To_Hex_String(AND_u64_u64_364_wire));
      --
    end process; 
    -- binary operator AND_u64_u64_364_inst
    process(mycount_351) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mycount_351, konst_363_wire_constant, tmp_var);
      AND_u64_u64_364_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u64_u64_386_inst flow-through 
    process(AND_u64_u64_386_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:AND_u64_u64_386_inst:flowthrough inputs: " & " nmycount_373 = "& Convert_SLV_To_Hex_String(nmycount_373) & " konst_385_wire_constant = "& Convert_SLV_To_Hex_String(konst_385_wire_constant) & " outputs:" & " AND_u64_u64_386_wire= "  & Convert_SLV_To_Hex_String(AND_u64_u64_386_wire));
      --
    end process; 
    -- binary operator AND_u64_u64_386_inst
    process(nmycount_373) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(nmycount_373, konst_385_wire_constant, tmp_var);
      AND_u64_u64_386_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u64_u1_342_inst flow-through 
    process(first_fill_343) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:EQ_u64_u1_342_inst:flowthrough inputs: " & " start_add_buffer = "& Convert_SLV_To_Hex_String(start_add_buffer) & " konst_341_wire_constant = "& Convert_SLV_To_Hex_String(konst_341_wire_constant) & " outputs:" & " first_fill_343= "  & Convert_SLV_To_Hex_String(first_fill_343));
      --
    end process; 
    -- binary operator EQ_u64_u1_342_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_341_wire_constant, tmp_var);
      first_fill_343 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u64_u1_388_inst flow-through 
    process(fn_389) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:EQ_u64_u1_388_inst:flowthrough inputs: " & " AND_u64_u64_386_wire = "& Convert_SLV_To_Hex_String(AND_u64_u64_386_wire) & " konst_387_wire_constant = "& Convert_SLV_To_Hex_String(konst_387_wire_constant) & " outputs:" & " fn_389= "  & Convert_SLV_To_Hex_String(fn_389));
      --
    end process; 
    -- binary operator EQ_u64_u1_388_inst
    process(AND_u64_u64_386_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(AND_u64_u64_386_wire, konst_387_wire_constant, tmp_var);
      fn_389 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u64_u64_326_inst flow-through 
    process(sh_start_327) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:LSHR_u64_u64_326_inst:flowthrough inputs: " & " start_add_buffer = "& Convert_SLV_To_Hex_String(start_add_buffer) & " konst_325_wire_constant = "& Convert_SLV_To_Hex_String(konst_325_wire_constant) & " outputs:" & " sh_start_327= "  & Convert_SLV_To_Hex_String(sh_start_327));
      --
    end process; 
    -- binary operator LSHR_u64_u64_326_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(start_add_buffer, konst_325_wire_constant, tmp_var);
      sh_start_327 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u64_u64_377_inst flow-through 
    process(LSHR_u64_u64_377_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:LSHR_u64_u64_377_inst:flowthrough inputs: " & " fetch_val_355 = "& Convert_SLV_To_Hex_String(fetch_val_355) & " my_num1_368 = "& Convert_SLV_To_Hex_String(my_num1_368) & " outputs:" & " LSHR_u64_u64_377_wire= "  & Convert_SLV_To_Hex_String(LSHR_u64_u64_377_wire));
      --
    end process; 
    -- binary operator LSHR_u64_u64_377_inst
    process(fetch_val_355, my_num1_368) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val_355, my_num1_368, tmp_var);
      LSHR_u64_u64_377_wire <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u64_u64_395_inst flow-through 
    process(LSHR_u64_u64_395_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:LSHR_u64_u64_395_inst:flowthrough inputs: " & " nmycount_373 = "& Convert_SLV_To_Hex_String(nmycount_373) & " konst_394_wire_constant = "& Convert_SLV_To_Hex_String(konst_394_wire_constant) & " outputs:" & " LSHR_u64_u64_395_wire= "  & Convert_SLV_To_Hex_String(LSHR_u64_u64_395_wire));
      --
    end process; 
    -- binary operator LSHR_u64_u64_395_inst
    process(nmycount_373) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nmycount_373, konst_394_wire_constant, tmp_var);
      LSHR_u64_u64_395_wire <= tmp_var; --
    end process;
    -- logger for split-operator SHL_u64_u64_367_inst flow-through 
    process(my_num1_368) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:SHL_u64_u64_367_inst:flowthrough inputs: " & " SUB_u64_u64_365_wire = "& Convert_SLV_To_Hex_String(SUB_u64_u64_365_wire) & " konst_366_wire_constant = "& Convert_SLV_To_Hex_String(konst_366_wire_constant) & " outputs:" & " my_num1_368= "  & Convert_SLV_To_Hex_String(my_num1_368));
      --
    end process; 
    -- binary operator SHL_u64_u64_367_inst
    process(SUB_u64_u64_365_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_365_wire, konst_366_wire_constant, tmp_var);
      my_num1_368 <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u64_u64_365_inst flow-through 
    process(SUB_u64_u64_365_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:SUB_u64_u64_365_inst:flowthrough inputs: " & " konst_361_wire_constant = "& Convert_SLV_To_Hex_String(konst_361_wire_constant) & " AND_u64_u64_364_wire = "& Convert_SLV_To_Hex_String(AND_u64_u64_364_wire) & " outputs:" & " SUB_u64_u64_365_wire= "  & Convert_SLV_To_Hex_String(SUB_u64_u64_365_wire));
      --
    end process; 
    -- binary operator SUB_u64_u64_365_inst
    process(konst_361_wire_constant, AND_u64_u64_364_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_361_wire_constant, AND_u64_u64_364_wire, tmp_var);
      SUB_u64_u64_365_wire <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u64_u64_423_inst flow-through 
    process(SUB_u64_u64_423_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:SUB_u64_u64_423_inst:flowthrough inputs: " & " end_add_buffer = "& Convert_SLV_To_Hex_String(end_add_buffer) & " konst_422_wire_constant = "& Convert_SLV_To_Hex_String(konst_422_wire_constant) & " outputs:" & " SUB_u64_u64_423_wire= "  & Convert_SLV_To_Hex_String(SUB_u64_u64_423_wire));
      --
    end process; 
    -- binary operator SUB_u64_u64_423_inst
    process(end_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, konst_422_wire_constant, tmp_var);
      SUB_u64_u64_423_wire <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u64_u64_430_inst flow-through 
    process(SUB_u64_u64_430_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:SUB_u64_u64_430_inst:flowthrough inputs: " & " first_fill_343 (guard)= " & Convert_SLV_To_String(first_fill_343) & " end_add_buffer = "& Convert_SLV_To_Hex_String(end_add_buffer) & " start_add_buffer = "& Convert_SLV_To_Hex_String(start_add_buffer) & " outputs:" & " SUB_u64_u64_430_wire= "  & Convert_SLV_To_Hex_String(SUB_u64_u64_430_wire));
      --
    end process; 
    -- binary operator SUB_u64_u64_430_inst
    process(end_add_buffer, start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, start_add_buffer, tmp_var);
      SUB_u64_u64_430_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u64_u1_424_inst flow-through 
    process(ULT_u64_u1_424_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ULT_u64_u1_424_inst:flowthrough inputs: " & " mycount_351 = "& Convert_SLV_To_Hex_String(mycount_351) & " SUB_u64_u64_423_wire = "& Convert_SLV_To_Hex_String(SUB_u64_u64_423_wire) & " outputs:" & " ULT_u64_u1_424_wire= "  & Convert_SLV_To_Hex_String(ULT_u64_u1_424_wire));
      --
    end process; 
    -- binary operator ULT_u64_u1_424_inst
    process(mycount_351, SUB_u64_u64_423_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_351, SUB_u64_u64_423_wire, tmp_var);
      ULT_u64_u1_424_wire <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_332_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_332_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:array_obj_ref_332_index_offset:started:   inputs: " & " R_sh_start_331_scaled = "& Convert_SLV_To_Hex_String(R_sh_start_331_scaled) & " array_obj_ref_332_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_332_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_332_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:array_obj_ref_332_index_offset:finished:  outputs: " & " array_obj_ref_332_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_332_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (13) : array_obj_ref_332_index_offset 
    ApIntAdd_group_13: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_sh_start_331_scaled;
      array_obj_ref_332_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_332_index_offset_req_0;
      array_obj_ref_332_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_332_index_offset_req_1;
      array_obj_ref_332_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_13_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- logger for split-operator array_obj_ref_396_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_396_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:array_obj_ref_396_index_offset:started:   inputs: " & " LSHR_u64_u64_395_scaled = "& Convert_SLV_To_Hex_String(LSHR_u64_u64_395_scaled) & " array_obj_ref_396_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_396_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_396_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:array_obj_ref_396_index_offset:finished:  outputs: " & " array_obj_ref_396_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_396_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (14) : array_obj_ref_396_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_395_scaled;
      array_obj_ref_396_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_396_index_offset_req_0;
      array_obj_ref_396_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_396_index_offset_req_1;
      array_obj_ref_396_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- logger for split-operator ptr_deref_337_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_337_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ptr_deref_337_load_0:started:   inputs: " & " ptr_deref_337_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_337_word_address_0));
          --
        end if; 
        if ptr_deref_337_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ptr_deref_337_load_0:finished:  outputs: " & " ptr_deref_337_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_337_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_405_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_405_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ptr_deref_405_load_0:started:   inputs: " & " fn_387_delayed_7_0_401 (guard)= " & Convert_SLV_To_String(fn_387_delayed_7_0_401) & " ptr_deref_405_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_405_word_address_0));
          --
        end if; 
        if ptr_deref_405_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:ptr_deref_405_load_0:finished:  outputs: " & " ptr_deref_405_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_405_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : ptr_deref_337_load_0 ptr_deref_405_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_337_load_0_req_0,
        ptr_deref_337_load_0_ack_0,
        ptr_deref_337_load_0_req_1,
        ptr_deref_337_load_0_ack_1,
        "ptr_deref_337_load_0",
        "memory_space_0" ,
        ptr_deref_337_data_0,
        ptr_deref_337_word_address_0,
        "ptr_deref_337_data_0",
        "ptr_deref_337_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_405_load_0_req_0,
        ptr_deref_405_load_0_ack_0,
        ptr_deref_405_load_0_req_1,
        ptr_deref_405_load_0_ack_1,
        "ptr_deref_405_load_0",
        "memory_space_0" ,
        ptr_deref_405_data_0,
        ptr_deref_405_word_address_0,
        "ptr_deref_405_data_0",
        "ptr_deref_405_word_address_0" -- 
      );
      reqL_unguarded(1) <= ptr_deref_337_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_405_load_0_req_0;
      ptr_deref_337_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_405_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_337_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_405_load_0_req_1;
      ptr_deref_337_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_405_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn_387_delayed_7_0_401(0);
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_337_word_address_0 & ptr_deref_405_word_address_0;
      ptr_deref_337_data_0 <= data_out(127 downto 64);
      ptr_deref_405_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator RPIPE_input_done_pipe_346_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_input_done_pipe_346_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:RPIPE_input_done_pipe_346_inst:started:   PipeRead from input_done_pipe inputs: " & " first_fill_343 (guard complement )= " & Convert_SLV_To_String(first_fill_343));
          --
        end if; 
        if RPIPE_input_done_pipe_346_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:RPIPE_input_done_pipe_346_inst:finished:  outputs: " & " start_next_347= "  & Convert_SLV_To_Hex_String(start_next_347));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_input_done_pipe_346_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_346_inst_req_0;
      RPIPE_input_done_pipe_346_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_346_inst_req_1;
      RPIPE_input_done_pipe_346_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_343(0);
      start_next_347 <= data_out(0 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_kernel_pipe1_380_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_kernel_pipe1_380_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:WPIPE_kernel_pipe1_380_inst:started:   PipeWrite to kernel_pipe1 inputs: " & " var_val_379 = "& Convert_SLV_To_Hex_String(var_val_379));
          --
        end if; 
        if WPIPE_kernel_pipe1_380_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:WPIPE_kernel_pipe1_380_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_380_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_380_inst_req_0;
      WPIPE_kernel_pipe1_380_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_380_inst_req_1;
      WPIPE_kernel_pipe1_380_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= var_val_379;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator WPIPE_size_pipe_427_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_size_pipe_427_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:WPIPE_size_pipe_427_inst:started:   PipeWrite to size_pipe inputs: " & " first_fill_343 (guard)= " & Convert_SLV_To_String(first_fill_343) & " type_cast_431_wire = "& Convert_SLV_To_Hex_String(type_cast_431_wire));
          --
        end if; 
        if WPIPE_size_pipe_427_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadKernelChannel:DP:WPIPE_size_pipe_427_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (1) : WPIPE_size_pipe_427_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_427_inst_req_0;
      WPIPE_size_pipe_427_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_427_inst_req_1;
      WPIPE_size_pipe_427_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= first_fill_343(0);
      data_in <= type_cast_431_wire;
      size_pipe_write_1_gI: SplitGuardInterface generic map(name => "size_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_637_start: Boolean;
  signal timer_CP_637_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_317_load_0_req_0 : boolean;
  signal LOAD_count_317_load_0_ack_0 : boolean;
  signal LOAD_count_317_load_0_req_1 : boolean;
  signal LOAD_count_317_load_0_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_637_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,timer_CP_637_start,"timer cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,timer_CP_637_symbol, "timer cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_637: Block -- control-path 
    signal timer_CP_637_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_637_elements(0) <= timer_CP_637_start;
    timer_CP_637_symbol <= timer_CP_637_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_318/$entry
      -- CP-element group 0: 	 assign_stmt_318/LOAD_count_317_sample_start_
      -- CP-element group 0: 	 assign_stmt_318/LOAD_count_317_update_start_
      -- CP-element group 0: 	 assign_stmt_318/LOAD_count_317_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_318/LOAD_count_317_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_318/LOAD_count_317_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_318/LOAD_count_317_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_318/LOAD_count_317_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_318/LOAD_count_317_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_318/LOAD_count_317_Update/$entry
      -- CP-element group 0: 	 assign_stmt_318/LOAD_count_317_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_318/LOAD_count_317_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_318/LOAD_count_317_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group timer_CP_637_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timer_CP_637_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:timer_CP_637_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:LOAD_count_317_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:LOAD_count_317_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => LOAD_count_317_load_0_req_1); -- 
    rr_658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => LOAD_count_317_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_318/LOAD_count_317_sample_completed_
      -- CP-element group 1: 	 assign_stmt_318/LOAD_count_317_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_318/LOAD_count_317_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_318/LOAD_count_317_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_318/LOAD_count_317_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group timer_CP_637_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timer_CP_637_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:timer_CP_637_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:LOAD_count_317_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_317_load_0_ack_0, ack => timer_CP_637_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_318/$exit
      -- CP-element group 2: 	 assign_stmt_318/LOAD_count_317_update_completed_
      -- CP-element group 2: 	 assign_stmt_318/LOAD_count_317_Update/$exit
      -- CP-element group 2: 	 assign_stmt_318/LOAD_count_317_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_318/LOAD_count_317_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_318/LOAD_count_317_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_318/LOAD_count_317_Update/LOAD_count_317_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_318/LOAD_count_317_Update/LOAD_count_317_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_318/LOAD_count_317_Update/LOAD_count_317_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_318/LOAD_count_317_Update/LOAD_count_317_Merge/merge_ack
      -- 
    -- logger for CP element group timer_CP_637_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timer_CP_637_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:timer_CP_637_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:LOAD_count_317_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_317_load_0_ack_1, ack => timer_CP_637_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_317_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_317_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_317_word_address_0 <= "0";
    -- logger for operator LOAD_count_317_gather_scatter flow-through 
    process(c_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:timer:DP:LOAD_count_317_gather_scatter:flowthrough  inputs: " & " LOAD_count_317_data_0 = "& Convert_SLV_To_Hex_String(LOAD_count_317_data_0) & "outputs: " & " c_buffer= "  & Convert_SLV_To_Hex_String(c_buffer));
      --
    end process; 
    -- equivalence LOAD_count_317_gather_scatter
    process(LOAD_count_317_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_317_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- logger for split-operator LOAD_count_317_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_count_317_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:timer:DP:LOAD_count_317_load_0:started:   inputs: " & " LOAD_count_317_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_count_317_word_address_0));
          --
        end if; 
        if LOAD_count_317_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:timer:DP:LOAD_count_317_load_0:finished:  outputs: " & " LOAD_count_317_data_0= "  & Convert_SLV_To_Hex_String(LOAD_count_317_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : LOAD_count_317_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_count_317_load_0_req_0,
        LOAD_count_317_load_0_ack_0,
        LOAD_count_317_load_0_req_1,
        LOAD_count_317_load_0_ack_1,
        "LOAD_count_317_load_0",
        "memory_space_2" ,
        LOAD_count_317_data_0,
        LOAD_count_317_word_address_0,
        "LOAD_count_317_data_0",
        "LOAD_count_317_word_address_0" -- 
      );
      reqL_unguarded(0) <= LOAD_count_317_load_0_req_0;
      LOAD_count_317_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_317_load_0_req_1;
      LOAD_count_317_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_317_word_address_0;
      LOAD_count_317_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_3899_start: Boolean;
  signal timerDaemon_CP_3899_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_1630_req_0 : boolean;
  signal do_while_stmt_1628_branch_ack_0 : boolean;
  signal ADD_u64_u64_1636_inst_ack_1 : boolean;
  signal do_while_stmt_1628_branch_req_0 : boolean;
  signal do_while_stmt_1628_branch_ack_1 : boolean;
  signal phi_stmt_1630_ack_0 : boolean;
  signal phi_stmt_1630_req_1 : boolean;
  signal ADD_u64_u64_1636_inst_req_1 : boolean;
  signal ADD_u64_u64_1636_inst_ack_0 : boolean;
  signal ADD_u64_u64_1636_inst_req_0 : boolean;
  signal STORE_count_1638_store_0_ack_1 : boolean;
  signal STORE_count_1638_store_0_req_1 : boolean;
  signal STORE_count_1638_store_0_ack_0 : boolean;
  signal STORE_count_1638_store_0_req_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_3899_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3899_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_3899_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3899_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,timerDaemon_CP_3899_start,"timerDaemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,timerDaemon_CP_3899_symbol, "timerDaemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_3899: Block -- control-path 
    signal timerDaemon_CP_3899_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_3899_elements(0) <= timerDaemon_CP_3899_start;
    timerDaemon_CP_3899_symbol <= timerDaemon_CP_3899_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1627/do_while_stmt_1628__entry__
      -- CP-element group 0: 	 branch_block_stmt_1627/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1627/branch_block_stmt_1627__entry__
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	39 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1627/do_while_stmt_1628__exit__
      -- CP-element group 1: 	 branch_block_stmt_1627/branch_block_stmt_1627__exit__
      -- CP-element group 1: 	 branch_block_stmt_1627/$exit
      -- CP-element group 1: 	 $exit
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_3899_elements(1) <= timerDaemon_CP_3899_elements(39);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628__entry__
      -- CP-element group 2: 	 branch_block_stmt_1627/do_while_stmt_1628/$entry
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_3899_elements(2) <= timerDaemon_CP_3899_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	39 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628__exit__
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_3899_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1627/do_while_stmt_1628/loop_back
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_3899_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	37 
    -- CP-element group 5: 	38 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1627/do_while_stmt_1628/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1627/do_while_stmt_1628/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1627/do_while_stmt_1628/loop_exit/$entry
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_3899_elements(5) <= timerDaemon_CP_3899_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	36 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1627/do_while_stmt_1628/loop_body_done
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_3899_elements(6) <= timerDaemon_CP_3899_elements(36);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_3899_elements(7) <= timerDaemon_CP_3899_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_3899_elements(8) <= timerDaemon_CP_3899_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	31 
    -- CP-element group 9: 	35 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_root_address_calculated
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_3899_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	35 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/condition_evaluated
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:do_while_stmt_1628_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3899_elements(10), ack => do_while_stmt_1628_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3899_elements(15) & timerDaemon_CP_3899_elements(35);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3899_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_sample_start__ps
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3899_elements(12) & timerDaemon_CP_3899_elements(15);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3899_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_sample_start_
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3899_elements(9) & timerDaemon_CP_3899_elements(14);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3899_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_update_start_
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3899_elements(9) & timerDaemon_CP_3899_elements(33);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3899_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_sample_completed__ps
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_3899_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	31 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_update_completed__ps
      -- CP-element group 15: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_update_completed_
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_3899_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_loopback_trigger
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_3899_elements(16) <= timerDaemon_CP_3899_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_loopback_sample_req_ps
      -- CP-element group 17: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_loopback_sample_req
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:phi_stmt_1630_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1630_loopback_sample_req_3938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1630_loopback_sample_req_3938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3899_elements(17), ack => phi_stmt_1630_req_1); -- 
    -- Element group timerDaemon_CP_3899_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_entry_trigger
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_3899_elements(18) <= timerDaemon_CP_3899_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_entry_sample_req_ps
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:phi_stmt_1630_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1630_entry_sample_req_3941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1630_entry_sample_req_3941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3899_elements(19), ack => phi_stmt_1630_req_0); -- 
    -- Element group timerDaemon_CP_3899_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_phi_mux_ack_ps
      -- CP-element group 20: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/phi_stmt_1630_phi_mux_ack
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:phi_stmt_1630_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1630_phi_mux_ack_3944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1630_ack_0, ack => timerDaemon_CP_3899_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/type_cast_1633_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/type_cast_1633_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/type_cast_1633_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/type_cast_1633_sample_start__ps
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_3899_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/type_cast_1633_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/type_cast_1633_update_start__ps
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(22) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_3899_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/type_cast_1633_update_completed__ps
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(23) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_3899_elements(23) <= timerDaemon_CP_3899_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/type_cast_1633_update_completed_
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_3899_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => timerDaemon_CP_3899_elements(22), ack => timerDaemon_CP_3899_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_sample_start__ps
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_3899_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_update_start__ps
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(26) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_3899_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_sample_start_
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:ADD_u64_u64_1636_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3899_elements(27), ack => ADD_u64_u64_1636_inst_req_0); -- 
    timerDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3899_elements(25) & timerDaemon_CP_3899_elements(29);
      gj_timerDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3899_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_update_start_
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:ADD_u64_u64_1636_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3899_elements(28), ack => ADD_u64_u64_1636_inst_req_1); -- 
    timerDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3899_elements(26) & timerDaemon_CP_3899_elements(30);
      gj_timerDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3899_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_sample_completed_
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:ADD_u64_u64_1636_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1636_inst_ack_0, ack => timerDaemon_CP_3899_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/ADD_u64_u64_1636_update_completed__ps
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:ADD_u64_u64_1636_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1636_inst_ack_1, ack => timerDaemon_CP_3899_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	15 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Sample/STORE_count_1638_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Sample/STORE_count_1638_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Sample/STORE_count_1638_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Sample/word_access_start/word_0/rr
      -- CP-element group 31: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Sample/STORE_count_1638_Split/split_ack
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:STORE_count_1638_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3899_elements(31), ack => STORE_count_1638_store_0_req_0); -- 
    timerDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_3899_elements(9) & timerDaemon_CP_3899_elements(15) & timerDaemon_CP_3899_elements(33);
      gj_timerDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3899_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Update/word_access_complete/word_0/cr
      -- CP-element group 32: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Update/$entry
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:STORE_count_1638_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3899_elements(32), ack => STORE_count_1638_store_0_req_1); -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= timerDaemon_CP_3899_elements(34);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3899_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Sample/word_access_start/word_0/ra
      -- CP-element group 33: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Sample/word_access_start/$exit
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:STORE_count_1638_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_1638_store_0_ack_0, ack => timerDaemon_CP_3899_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Update/word_access_complete/word_0/ca
      -- CP-element group 34: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/STORE_count_1638_Update/$exit
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:STORE_count_1638_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_1638_store_0_ack_1, ack => timerDaemon_CP_3899_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(35) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_3899_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => timerDaemon_CP_3899_elements(9), ack => timerDaemon_CP_3899_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	6 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1627/do_while_stmt_1628/do_while_stmt_1628_loop_body/$exit
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(36) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3899_elements(14) & timerDaemon_CP_3899_elements(34);
      gj_timerDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3899_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	5 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_1627/do_while_stmt_1628/loop_exit/$exit
      -- CP-element group 37: 	 branch_block_stmt_1627/do_while_stmt_1628/loop_exit/ack
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:do_while_stmt_1628_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1628_branch_ack_0, ack => timerDaemon_CP_3899_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_1627/do_while_stmt_1628/loop_taken/$exit
      -- CP-element group 38: 	 branch_block_stmt_1627/do_while_stmt_1628/loop_taken/ack
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:do_while_stmt_1628_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1628_branch_ack_1, ack => timerDaemon_CP_3899_elements(38)); -- 
    -- CP-element group 39:  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	3 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	1 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1627/do_while_stmt_1628/$exit
      -- 
    -- logger for CP element group timerDaemon_CP_3899_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_3899_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_3899_elements(39) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_3899_elements(39) <= timerDaemon_CP_3899_elements(3);
    timerDaemon_do_while_stmt_1628_terminator_4015: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_1628_terminator_4015", max_iterations_in_flight =>3) 
      port map(loop_body_exit => timerDaemon_CP_3899_elements(6),loop_continue => timerDaemon_CP_3899_elements(38),loop_terminate => timerDaemon_CP_3899_elements(37),loop_back => timerDaemon_CP_3899_elements(4),loop_exit => timerDaemon_CP_3899_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1630_phi_seq_3972_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_3899_elements(18);
      timerDaemon_CP_3899_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_3899_elements(21);
      timerDaemon_CP_3899_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_3899_elements(23);
      timerDaemon_CP_3899_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_3899_elements(16);
      timerDaemon_CP_3899_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_3899_elements(29);
      timerDaemon_CP_3899_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_3899_elements(30);
      timerDaemon_CP_3899_elements(17) <= phi_mux_reqs(1);
      phi_stmt_1630_phi_seq_3972 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_1630_phi_seq_3972") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_3899_elements(11), 
          phi_sample_ack => timerDaemon_CP_3899_elements(14), 
          phi_update_req => timerDaemon_CP_3899_elements(13), 
          phi_update_ack => timerDaemon_CP_3899_elements(15), 
          phi_mux_ack => timerDaemon_CP_3899_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3924_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_3899_elements(7);
        preds(1)  <= timerDaemon_CP_3899_elements(8);
        entry_tmerge_3924 : transition_merge -- 
          generic map(name => " entry_tmerge_3924")
          port map (preds => preds, symbol_out => timerDaemon_CP_3899_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u64_u64_1636_wire : std_logic_vector(63 downto 0);
    signal STORE_count_1638_data_0 : std_logic_vector(63 downto 0);
    signal STORE_count_1638_word_address_0 : std_logic_vector(0 downto 0);
    signal konst_1635_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1642_wire_constant : std_logic_vector(0 downto 0);
    signal ncount_1630 : std_logic_vector(63 downto 0);
    signal type_cast_1633_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_count_1638_word_address_0 <= "0";
    konst_1635_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_1642_wire_constant <= "1";
    type_cast_1633_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- logger for phi phi_stmt_1630
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1630_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:timerDaemon:DP:phi_stmt_1630:input-0 type_cast_1633_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1633_wire_constant));
          --
        end if;
        if phi_stmt_1630_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:timerDaemon:DP:phi_stmt_1630:input-1 ADD_u64_u64_1636_wire= " & Convert_SLV_To_Hex_String(ADD_u64_u64_1636_wire));
          --
        end if;
        if phi_stmt_1630_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:timerDaemon:DP:phi_stmt_1630:sample-completed");
          --
        end if;
        if phi_stmt_1630_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:timerDaemon:DP:phi_stmt_1630:output ncount_1630= " & Convert_SLV_To_Hex_String(ncount_1630));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1630: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1633_wire_constant & ADD_u64_u64_1636_wire;
      req <= phi_stmt_1630_req_0 & phi_stmt_1630_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1630",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1630_ack_0,
          idata => idata,
          odata => ncount_1630,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1630
    -- logger for operator STORE_count_1638_gather_scatter flow-through 
    process(STORE_count_1638_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:timerDaemon:DP:STORE_count_1638_gather_scatter:flowthrough  inputs: " & " ncount_1630 = "& Convert_SLV_To_Hex_String(ncount_1630) & "outputs: " & " STORE_count_1638_data_0= "  & Convert_SLV_To_Hex_String(STORE_count_1638_data_0));
      --
    end process; 
    -- equivalence STORE_count_1638_gather_scatter
    process(ncount_1630) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ncount_1630;
      ov(63 downto 0) := iv;
      STORE_count_1638_data_0 <= ov(63 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1628_branch_req_0," req0 do_while_stmt_1628_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1628_branch_ack_0," ack0 do_while_stmt_1628_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1628_branch_ack_1," ack1 do_while_stmt_1628_branch");
    do_while_stmt_1628_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1642_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1628_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1628_branch_req_0,
          ack0 => do_while_stmt_1628_branch_ack_0,
          ack1 => do_while_stmt_1628_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u64_u64_1636_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u64_u64_1636_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:timerDaemon:DP:ADD_u64_u64_1636_inst:started:   inputs: " & " ncount_1630 = "& Convert_SLV_To_Hex_String(ncount_1630) & " konst_1635_wire_constant = "& Convert_SLV_To_Hex_String(konst_1635_wire_constant));
          --
        end if; 
        if ADD_u64_u64_1636_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:timerDaemon:DP:ADD_u64_u64_1636_inst:finished:  outputs: " & " ADD_u64_u64_1636_wire= "  & Convert_SLV_To_Hex_String(ADD_u64_u64_1636_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : ADD_u64_u64_1636_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ncount_1630;
      ADD_u64_u64_1636_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1636_inst_req_0;
      ADD_u64_u64_1636_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1636_inst_req_1;
      ADD_u64_u64_1636_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator STORE_count_1638_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if STORE_count_1638_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:timerDaemon:DP:STORE_count_1638_store_0:started:   inputs: " & " STORE_count_1638_word_address_0 = "& Convert_SLV_To_Hex_String(STORE_count_1638_word_address_0) & " STORE_count_1638_data_0 = "& Convert_SLV_To_Hex_String(STORE_count_1638_data_0));
          --
        end if; 
        if STORE_count_1638_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:timerDaemon:DP:STORE_count_1638_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      STORE_count_1638_store_0_req_0,
      STORE_count_1638_store_0_ack_0,
      STORE_count_1638_store_0_req_1,
      STORE_count_1638_store_0_ack_1,
      "STORE_count_1638_store_0",
      "memory_space_2" ,
      STORE_count_1638_data_0,
      STORE_count_1638_word_address_0,
      "STORE_count_1638_data_0",
      "STORE_count_1638_word_address_0" -- 
    );
    -- shared store operator group (0) : STORE_count_1638_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_count_1638_store_0_req_0;
      STORE_count_1638_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_count_1638_store_0_req_1;
      STORE_count_1638_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_count_1638_word_address_0;
      data_in <= STORE_count_1638_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(15 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(15 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_num_cont :  std_logic_vector(15 downto 0);
  signal access_T_row1 :  std_logic_vector(15 downto 0);
  signal access_T_col1 :  std_logic_vector(15 downto 0);
  signal access_T_rk1 :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(95 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(95 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(95 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(127 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_end_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(127 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(127 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(31 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(1 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_num_cont <= access_T_in_args(95 downto 80);
  access_T_row1 <= access_T_in_args(79 downto 64);
  access_T_col1 <= access_T_in_args(63 downto 48);
  access_T_rk1 <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 96,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      num_cont => access_T_num_cont,
      row1 => access_T_row1,
      col1 => access_T_col1,
      rk1 => access_T_rk1,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(15 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(15 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(31 downto 16),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(95 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(127 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(15 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(31 downto 0),
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(15 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(0 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(15 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(127 downto 64);
  loadKernelChannel_end_add <= loadKernelChannel_in_args(63 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 128,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      end_add => loadKernelChannel_end_add,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(0 downto 0),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(31 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(1 downto 1),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(1 downto 1),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(31 downto 16),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
