-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_data : in   std_logic_vector(15 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_3522_start: Boolean;
  signal convTranspose_CP_3522_symbol: Boolean;
  -- volatile/operator module components. 
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_Block1_start_1208_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1208_inst_ack_1 : boolean;
  signal call_stmt_1203_call_req_0 : boolean;
  signal call_stmt_1203_call_ack_0 : boolean;
  signal WPIPE_Block1_start_1208_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1208_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1205_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1205_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1205_inst_req_1 : boolean;
  signal call_stmt_1203_call_req_1 : boolean;
  signal call_stmt_1203_call_ack_1 : boolean;
  signal WPIPE_Block0_start_1205_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1211_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1211_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1211_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1211_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1214_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1214_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1214_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1214_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1218_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1218_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1218_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1218_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1221_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1221_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1221_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1221_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1224_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1224_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1224_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1224_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1227_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1227_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1227_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1227_inst_ack_1 : boolean;
  signal call_stmt_1230_call_req_0 : boolean;
  signal call_stmt_1230_call_ack_0 : boolean;
  signal call_stmt_1230_call_req_1 : boolean;
  signal call_stmt_1230_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_3522_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3522_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_3522_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3522_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_3522: Block -- control-path 
    signal convTranspose_CP_3522_elements: BooleanArray(21 downto 0);
    -- 
  begin -- 
    convTranspose_CP_3522_elements(0) <= convTranspose_CP_3522_start;
    convTranspose_CP_3522_symbol <= convTranspose_CP_3522_elements(21);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_1201/call_stmt_1203/$entry
      -- CP-element group 0: 	 branch_block_stmt_1201/$entry
      -- CP-element group 0: 	 branch_block_stmt_1201/branch_block_stmt_1201__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1201/call_stmt_1203/call_stmt_1203_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1201/call_stmt_1203/call_stmt_1203_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1201/call_stmt_1203/call_stmt_1203_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_1201/call_stmt_1203__entry__
      -- CP-element group 0: 	 branch_block_stmt_1201/call_stmt_1203/call_stmt_1203_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1201/call_stmt_1203/call_stmt_1203_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1201/call_stmt_1203/call_stmt_1203_Update/ccr
      -- 
    crr_3548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(0), ack => call_stmt_1203_call_req_0); -- 
    ccr_3553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(0), ack => call_stmt_1203_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_1201/call_stmt_1203/call_stmt_1203_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1201/call_stmt_1203/call_stmt_1203_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1201/call_stmt_1203/call_stmt_1203_Sample/cra
      -- 
    cra_3549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1203_call_ack_0, ack => convTranspose_CP_3522_elements(1)); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	13 
    -- CP-element group 2:  members (31) 
      -- CP-element group 2: 	 branch_block_stmt_1201/call_stmt_1203/$exit
      -- CP-element group 2: 	 branch_block_stmt_1201/call_stmt_1203/call_stmt_1203_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1201/call_stmt_1203__exit__
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block1_start_1208_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block0_start_1205_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block1_start_1208_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block1_start_1208_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1201/call_stmt_1203/call_stmt_1203_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block0_start_1205_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block0_start_1205_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block2_start_1211_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1201/call_stmt_1203/call_stmt_1203_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/$entry
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228__entry__
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block2_start_1211_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block2_start_1211_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block3_start_1214_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block3_start_1214_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block3_start_1214_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block0_done_1218_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block0_done_1218_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block0_done_1218_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block1_done_1221_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block1_done_1221_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block1_done_1221_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block2_done_1224_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block2_done_1224_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block2_done_1224_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block3_done_1227_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block3_done_1227_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block3_done_1227_Sample/rr
      -- 
    cca_3554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1203_call_ack_1, ack => convTranspose_CP_3522_elements(2)); -- 
    req_3579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(2), ack => WPIPE_Block1_start_1208_inst_req_0); -- 
    req_3565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(2), ack => WPIPE_Block0_start_1205_inst_req_0); -- 
    req_3593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(2), ack => WPIPE_Block2_start_1211_inst_req_0); -- 
    req_3607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(2), ack => WPIPE_Block3_start_1214_inst_req_0); -- 
    rr_3621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(2), ack => RPIPE_Block0_done_1218_inst_req_0); -- 
    rr_3635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(2), ack => RPIPE_Block1_done_1221_inst_req_0); -- 
    rr_3649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(2), ack => RPIPE_Block2_done_1224_inst_req_0); -- 
    rr_3663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(2), ack => RPIPE_Block3_done_1227_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block0_start_1205_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block0_start_1205_Sample/ack
      -- CP-element group 3: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block0_start_1205_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block0_start_1205_Update/req
      -- CP-element group 3: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block0_start_1205_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block0_start_1205_update_start_
      -- 
    ack_3566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1205_inst_ack_0, ack => convTranspose_CP_3522_elements(3)); -- 
    req_3570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(3), ack => WPIPE_Block0_start_1205_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	19 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block0_start_1205_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block0_start_1205_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block0_start_1205_Update/ack
      -- 
    ack_3571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1205_inst_ack_1, ack => convTranspose_CP_3522_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block1_start_1208_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block1_start_1208_Update/req
      -- CP-element group 5: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block1_start_1208_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block1_start_1208_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block1_start_1208_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block1_start_1208_Sample/ack
      -- 
    ack_3580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1208_inst_ack_0, ack => convTranspose_CP_3522_elements(5)); -- 
    req_3584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(5), ack => WPIPE_Block1_start_1208_inst_req_1); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	19 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block1_start_1208_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block1_start_1208_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block1_start_1208_update_completed_
      -- 
    ack_3585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1208_inst_ack_1, ack => convTranspose_CP_3522_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block2_start_1211_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block2_start_1211_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block2_start_1211_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block2_start_1211_Sample/ack
      -- CP-element group 7: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block2_start_1211_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block2_start_1211_Update/req
      -- 
    ack_3594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1211_inst_ack_0, ack => convTranspose_CP_3522_elements(7)); -- 
    req_3598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(7), ack => WPIPE_Block2_start_1211_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	19 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block2_start_1211_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block2_start_1211_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block2_start_1211_Update/ack
      -- 
    ack_3599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1211_inst_ack_1, ack => convTranspose_CP_3522_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block3_start_1214_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block3_start_1214_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block3_start_1214_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block3_start_1214_Sample/ack
      -- CP-element group 9: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block3_start_1214_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block3_start_1214_Update/req
      -- 
    ack_3608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1214_inst_ack_0, ack => convTranspose_CP_3522_elements(9)); -- 
    req_3612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(9), ack => WPIPE_Block3_start_1214_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	19 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block3_start_1214_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block3_start_1214_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/WPIPE_Block3_start_1214_Update/ack
      -- 
    ack_3613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1214_inst_ack_1, ack => convTranspose_CP_3522_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block0_done_1218_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block0_done_1218_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block0_done_1218_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block0_done_1218_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block0_done_1218_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block0_done_1218_Update/cr
      -- 
    ra_3622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1218_inst_ack_0, ack => convTranspose_CP_3522_elements(11)); -- 
    cr_3626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(11), ack => RPIPE_Block0_done_1218_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	19 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block0_done_1218_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block0_done_1218_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block0_done_1218_Update/ca
      -- 
    ca_3627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1218_inst_ack_1, ack => convTranspose_CP_3522_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block1_done_1221_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block1_done_1221_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block1_done_1221_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block1_done_1221_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block1_done_1221_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block1_done_1221_Update/cr
      -- 
    ra_3636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1221_inst_ack_0, ack => convTranspose_CP_3522_elements(13)); -- 
    cr_3640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(13), ack => RPIPE_Block1_done_1221_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	19 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block1_done_1221_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block1_done_1221_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block1_done_1221_Update/ca
      -- 
    ca_3641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1221_inst_ack_1, ack => convTranspose_CP_3522_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block2_done_1224_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block2_done_1224_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block2_done_1224_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block2_done_1224_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block2_done_1224_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block2_done_1224_Update/cr
      -- 
    ra_3650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1224_inst_ack_0, ack => convTranspose_CP_3522_elements(15)); -- 
    cr_3654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(15), ack => RPIPE_Block2_done_1224_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	19 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block2_done_1224_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block2_done_1224_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block2_done_1224_Update/ca
      -- 
    ca_3655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1224_inst_ack_1, ack => convTranspose_CP_3522_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block3_done_1227_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block3_done_1227_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block3_done_1227_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block3_done_1227_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block3_done_1227_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block3_done_1227_Update/cr
      -- 
    ra_3664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1227_inst_ack_0, ack => convTranspose_CP_3522_elements(17)); -- 
    cr_3668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(17), ack => RPIPE_Block3_done_1227_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block3_done_1227_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block3_done_1227_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/RPIPE_Block3_done_1227_Update/ca
      -- 
    ca_3669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1227_inst_ack_1, ack => convTranspose_CP_3522_elements(18)); -- 
    -- CP-element group 19:  join  fork  transition  place  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	6 
    -- CP-element group 19: 	10 
    -- CP-element group 19: 	14 
    -- CP-element group 19: 	4 
    -- CP-element group 19: 	8 
    -- CP-element group 19: 	12 
    -- CP-element group 19: 	18 
    -- CP-element group 19: 	16 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (10) 
      -- CP-element group 19: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228__exit__
      -- CP-element group 19: 	 branch_block_stmt_1201/call_stmt_1230__entry__
      -- CP-element group 19: 	 branch_block_stmt_1201/assign_stmt_1207_to_assign_stmt_1228/$exit
      -- CP-element group 19: 	 branch_block_stmt_1201/call_stmt_1230/$entry
      -- CP-element group 19: 	 branch_block_stmt_1201/call_stmt_1230/call_stmt_1230_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1201/call_stmt_1230/call_stmt_1230_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1201/call_stmt_1230/call_stmt_1230_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1201/call_stmt_1230/call_stmt_1230_Sample/crr
      -- CP-element group 19: 	 branch_block_stmt_1201/call_stmt_1230/call_stmt_1230_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1201/call_stmt_1230/call_stmt_1230_Update/ccr
      -- 
    crr_3680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(19), ack => call_stmt_1230_call_req_0); -- 
    ccr_3685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3522_elements(19), ack => call_stmt_1230_call_req_1); -- 
    convTranspose_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= convTranspose_CP_3522_elements(6) & convTranspose_CP_3522_elements(10) & convTranspose_CP_3522_elements(14) & convTranspose_CP_3522_elements(4) & convTranspose_CP_3522_elements(8) & convTranspose_CP_3522_elements(12) & convTranspose_CP_3522_elements(18) & convTranspose_CP_3522_elements(16);
      gj_convTranspose_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_3522_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1201/call_stmt_1230/call_stmt_1230_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1201/call_stmt_1230/call_stmt_1230_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1201/call_stmt_1230/call_stmt_1230_Sample/cra
      -- 
    cra_3681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1230_call_ack_0, ack => convTranspose_CP_3522_elements(20)); -- 
    -- CP-element group 21:  transition  place  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (16) 
      -- CP-element group 21: 	 branch_block_stmt_1201/$exit
      -- CP-element group 21: 	 branch_block_stmt_1201/merge_stmt_1232__exit__
      -- CP-element group 21: 	 branch_block_stmt_1201/branch_block_stmt_1201__exit__
      -- CP-element group 21: 	 $exit
      -- CP-element group 21: 	 branch_block_stmt_1201/call_stmt_1230__exit__
      -- CP-element group 21: 	 branch_block_stmt_1201/return__
      -- CP-element group 21: 	 branch_block_stmt_1201/call_stmt_1230/$exit
      -- CP-element group 21: 	 branch_block_stmt_1201/call_stmt_1230/call_stmt_1230_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1201/call_stmt_1230/call_stmt_1230_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1201/call_stmt_1230/call_stmt_1230_Update/cca
      -- CP-element group 21: 	 branch_block_stmt_1201/return___PhiReq/$entry
      -- CP-element group 21: 	 branch_block_stmt_1201/return___PhiReq/$exit
      -- CP-element group 21: 	 branch_block_stmt_1201/merge_stmt_1232_PhiReqMerge
      -- CP-element group 21: 	 branch_block_stmt_1201/merge_stmt_1232_PhiAck/$entry
      -- CP-element group 21: 	 branch_block_stmt_1201/merge_stmt_1232_PhiAck/$exit
      -- CP-element group 21: 	 branch_block_stmt_1201/merge_stmt_1232_PhiAck/dummy
      -- 
    cca_3686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1230_call_ack_1, ack => convTranspose_CP_3522_elements(21)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal call11_1228 : std_logic_vector(15 downto 0);
    signal call5_1219 : std_logic_vector(15 downto 0);
    signal call7_1222 : std_logic_vector(15 downto 0);
    signal call9_1225 : std_logic_vector(15 downto 0);
    signal call_1203 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    -- shared inport operator group (0) : RPIPE_Block0_done_1218_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1218_inst_req_0;
      RPIPE_Block0_done_1218_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1218_inst_req_1;
      RPIPE_Block0_done_1218_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call5_1219 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1221_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1221_inst_req_0;
      RPIPE_Block1_done_1221_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1221_inst_req_1;
      RPIPE_Block1_done_1221_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call7_1222 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1224_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1224_inst_req_0;
      RPIPE_Block2_done_1224_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1224_inst_req_1;
      RPIPE_Block2_done_1224_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call9_1225 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1227_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1227_inst_req_0;
      RPIPE_Block3_done_1227_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1227_inst_req_1;
      RPIPE_Block3_done_1227_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call11_1228 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_Block0_start_1205_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_start_1205_inst_req_0;
      WPIPE_Block0_start_1205_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_start_1205_inst_req_1;
      WPIPE_Block0_start_1205_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1203;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1208_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_start_1208_inst_req_0;
      WPIPE_Block1_start_1208_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_start_1208_inst_req_1;
      WPIPE_Block1_start_1208_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1203;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1211_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_start_1211_inst_req_0;
      WPIPE_Block2_start_1211_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_start_1211_inst_req_1;
      WPIPE_Block2_start_1211_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1203;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1214_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_start_1214_inst_req_0;
      WPIPE_Block3_start_1214_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_start_1214_inst_req_1;
      WPIPE_Block3_start_1214_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1203;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared call operator group (0) : call_stmt_1203_call 
    testConfigure_call_group_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1203_call_req_0;
      call_stmt_1203_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1203_call_req_1;
      call_stmt_1203_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_0_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_1203 <= data_out(15 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          dataL => testConfigure_return_data(15 downto 0),
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1230_call 
    sendOutput_call_group_1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1230_call_req_0;
      call_stmt_1230_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1230_call_req_1;
      call_stmt_1230_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_1_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3695_start: Boolean;
  signal convTransposeA_CP_3695_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1310_inst_req_1 : boolean;
  signal type_cast_1310_inst_ack_1 : boolean;
  signal ptr_deref_1322_load_0_req_0 : boolean;
  signal type_cast_1296_inst_ack_1 : boolean;
  signal ptr_deref_1289_load_0_ack_0 : boolean;
  signal ptr_deref_1263_load_0_ack_1 : boolean;
  signal ptr_deref_1346_load_0_ack_0 : boolean;
  signal ptr_deref_1306_load_0_req_1 : boolean;
  signal LOAD_padding_1292_load_0_req_0 : boolean;
  signal type_cast_1277_inst_req_0 : boolean;
  signal type_cast_1277_inst_ack_0 : boolean;
  signal type_cast_1277_inst_ack_1 : boolean;
  signal ptr_deref_1306_load_0_ack_1 : boolean;
  signal LOAD_padding_1292_load_0_ack_0 : boolean;
  signal ptr_deref_1334_load_0_ack_0 : boolean;
  signal ptr_deref_1346_load_0_ack_1 : boolean;
  signal ptr_deref_1334_load_0_req_0 : boolean;
  signal ptr_deref_1322_load_0_ack_0 : boolean;
  signal ptr_deref_1289_load_0_req_0 : boolean;
  signal type_cast_1296_inst_req_1 : boolean;
  signal type_cast_1277_inst_req_1 : boolean;
  signal ptr_deref_1263_load_0_req_0 : boolean;
  signal ptr_deref_1346_load_0_req_1 : boolean;
  signal type_cast_1296_inst_req_0 : boolean;
  signal ptr_deref_1263_load_0_req_1 : boolean;
  signal ptr_deref_1346_load_0_req_0 : boolean;
  signal ptr_deref_1263_load_0_ack_0 : boolean;
  signal type_cast_1296_inst_ack_0 : boolean;
  signal ptr_deref_1334_load_0_req_1 : boolean;
  signal ptr_deref_1334_load_0_ack_1 : boolean;
  signal type_cast_1310_inst_req_0 : boolean;
  signal ptr_deref_1289_load_0_req_1 : boolean;
  signal ptr_deref_1289_load_0_ack_1 : boolean;
  signal ptr_deref_1306_load_0_ack_0 : boolean;
  signal ptr_deref_1306_load_0_req_0 : boolean;
  signal ptr_deref_1273_load_0_ack_1 : boolean;
  signal ptr_deref_1273_load_0_req_1 : boolean;
  signal LOAD_padding_1292_load_0_ack_1 : boolean;
  signal LOAD_padding_1292_load_0_req_1 : boolean;
  signal ptr_deref_1322_load_0_ack_1 : boolean;
  signal ptr_deref_1322_load_0_req_1 : boolean;
  signal type_cast_1310_inst_ack_0 : boolean;
  signal ptr_deref_1273_load_0_ack_0 : boolean;
  signal ptr_deref_1273_load_0_req_0 : boolean;
  signal RPIPE_Block0_start_1238_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1238_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1238_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1238_inst_ack_1 : boolean;
  signal ptr_deref_1251_load_0_req_0 : boolean;
  signal ptr_deref_1251_load_0_ack_0 : boolean;
  signal ptr_deref_1251_load_0_req_1 : boolean;
  signal ptr_deref_1251_load_0_ack_1 : boolean;
  signal ptr_deref_1364_load_0_req_0 : boolean;
  signal ptr_deref_1364_load_0_ack_0 : boolean;
  signal ptr_deref_1364_load_0_req_1 : boolean;
  signal ptr_deref_1364_load_0_ack_1 : boolean;
  signal type_cast_1393_inst_req_0 : boolean;
  signal type_cast_1393_inst_ack_0 : boolean;
  signal type_cast_1393_inst_req_1 : boolean;
  signal type_cast_1393_inst_ack_1 : boolean;
  signal type_cast_1398_inst_req_0 : boolean;
  signal type_cast_1398_inst_ack_0 : boolean;
  signal type_cast_1398_inst_req_1 : boolean;
  signal type_cast_1398_inst_ack_1 : boolean;
  signal type_cast_1520_inst_req_0 : boolean;
  signal type_cast_1520_inst_ack_0 : boolean;
  signal type_cast_1520_inst_req_1 : boolean;
  signal type_cast_1520_inst_ack_1 : boolean;
  signal type_cast_1551_inst_req_0 : boolean;
  signal type_cast_1551_inst_ack_0 : boolean;
  signal type_cast_1551_inst_req_1 : boolean;
  signal type_cast_1551_inst_ack_1 : boolean;
  signal array_obj_ref_1557_index_offset_req_0 : boolean;
  signal array_obj_ref_1557_index_offset_ack_0 : boolean;
  signal array_obj_ref_1557_index_offset_req_1 : boolean;
  signal array_obj_ref_1557_index_offset_ack_1 : boolean;
  signal addr_of_1558_final_reg_req_0 : boolean;
  signal addr_of_1558_final_reg_ack_0 : boolean;
  signal addr_of_1558_final_reg_req_1 : boolean;
  signal addr_of_1558_final_reg_ack_1 : boolean;
  signal ptr_deref_1562_load_0_req_0 : boolean;
  signal ptr_deref_1562_load_0_ack_0 : boolean;
  signal ptr_deref_1562_load_0_req_1 : boolean;
  signal ptr_deref_1562_load_0_ack_1 : boolean;
  signal type_cast_1582_inst_req_0 : boolean;
  signal type_cast_1582_inst_ack_0 : boolean;
  signal type_cast_1582_inst_req_1 : boolean;
  signal type_cast_1582_inst_ack_1 : boolean;
  signal array_obj_ref_1588_index_offset_req_0 : boolean;
  signal array_obj_ref_1588_index_offset_ack_0 : boolean;
  signal array_obj_ref_1588_index_offset_req_1 : boolean;
  signal array_obj_ref_1588_index_offset_ack_1 : boolean;
  signal addr_of_1589_final_reg_req_0 : boolean;
  signal addr_of_1589_final_reg_ack_0 : boolean;
  signal addr_of_1589_final_reg_req_1 : boolean;
  signal addr_of_1589_final_reg_ack_1 : boolean;
  signal ptr_deref_1592_store_0_req_0 : boolean;
  signal ptr_deref_1592_store_0_ack_0 : boolean;
  signal ptr_deref_1592_store_0_req_1 : boolean;
  signal ptr_deref_1592_store_0_ack_1 : boolean;
  signal type_cast_1598_inst_req_0 : boolean;
  signal type_cast_1598_inst_ack_0 : boolean;
  signal type_cast_1598_inst_req_1 : boolean;
  signal type_cast_1598_inst_ack_1 : boolean;
  signal if_stmt_1611_branch_req_0 : boolean;
  signal if_stmt_1611_branch_ack_1 : boolean;
  signal if_stmt_1611_branch_ack_0 : boolean;
  signal type_cast_1635_inst_req_0 : boolean;
  signal type_cast_1635_inst_ack_0 : boolean;
  signal type_cast_1635_inst_req_1 : boolean;
  signal type_cast_1635_inst_ack_1 : boolean;
  signal type_cast_1644_inst_req_0 : boolean;
  signal type_cast_1644_inst_ack_0 : boolean;
  signal type_cast_1644_inst_req_1 : boolean;
  signal type_cast_1644_inst_ack_1 : boolean;
  signal type_cast_1661_inst_req_0 : boolean;
  signal type_cast_1661_inst_ack_0 : boolean;
  signal type_cast_1661_inst_req_1 : boolean;
  signal type_cast_1661_inst_ack_1 : boolean;
  signal if_stmt_1668_branch_req_0 : boolean;
  signal if_stmt_1668_branch_ack_1 : boolean;
  signal if_stmt_1668_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1676_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1676_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1676_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1676_inst_ack_1 : boolean;
  signal phi_stmt_1374_req_0 : boolean;
  signal phi_stmt_1381_req_0 : boolean;
  signal type_cast_1380_inst_req_0 : boolean;
  signal type_cast_1380_inst_ack_0 : boolean;
  signal type_cast_1380_inst_req_1 : boolean;
  signal type_cast_1380_inst_ack_1 : boolean;
  signal phi_stmt_1374_req_1 : boolean;
  signal type_cast_1387_inst_req_0 : boolean;
  signal type_cast_1387_inst_ack_0 : boolean;
  signal type_cast_1387_inst_req_1 : boolean;
  signal type_cast_1387_inst_ack_1 : boolean;
  signal phi_stmt_1381_req_1 : boolean;
  signal phi_stmt_1374_ack_0 : boolean;
  signal phi_stmt_1381_ack_0 : boolean;
  signal type_cast_1510_inst_req_0 : boolean;
  signal type_cast_1510_inst_ack_0 : boolean;
  signal type_cast_1510_inst_req_1 : boolean;
  signal type_cast_1510_inst_ack_1 : boolean;
  signal phi_stmt_1504_req_1 : boolean;
  signal phi_stmt_1504_req_0 : boolean;
  signal phi_stmt_1504_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3695_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3695_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3695_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3695_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3695: Block -- control-path 
    signal convTransposeA_CP_3695_elements: BooleanArray(88 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3695_elements(0) <= convTransposeA_CP_3695_start;
    convTransposeA_CP_3695_symbol <= convTransposeA_CP_3695_elements(68);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1236/$entry
      -- CP-element group 0: 	 branch_block_stmt_1236/branch_block_stmt_1236__entry__
      -- CP-element group 0: 	 branch_block_stmt_1236/assign_stmt_1239__entry__
      -- CP-element group 0: 	 branch_block_stmt_1236/assign_stmt_1239/$entry
      -- CP-element group 0: 	 branch_block_stmt_1236/assign_stmt_1239/RPIPE_Block0_start_1238_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1236/assign_stmt_1239/RPIPE_Block0_start_1238_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1236/assign_stmt_1239/RPIPE_Block0_start_1238_Sample/rr
      -- 
    rr_3743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(0), ack => RPIPE_Block0_start_1238_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1236/assign_stmt_1239/RPIPE_Block0_start_1238_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1236/assign_stmt_1239/RPIPE_Block0_start_1238_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1236/assign_stmt_1239/RPIPE_Block0_start_1238_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1236/assign_stmt_1239/RPIPE_Block0_start_1238_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1236/assign_stmt_1239/RPIPE_Block0_start_1238_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1236/assign_stmt_1239/RPIPE_Block0_start_1238_Update/cr
      -- 
    ra_3744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1238_inst_ack_0, ack => convTransposeA_CP_3695_elements(1)); -- 
    cr_3748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(1), ack => RPIPE_Block0_start_1238_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	16 
    -- CP-element group 2:  members (262) 
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1310_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1277_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1310_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1310_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1296_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1277_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1296_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1277_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1296_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1239__exit__
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371__entry__
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1239/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1239/RPIPE_Block0_start_1238_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1239/RPIPE_Block0_start_1238_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1239/RPIPE_Block0_start_1238_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Update/word_access_complete/word_0/cr
      -- 
    ca_3749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1238_inst_ack_1, ack => convTransposeA_CP_3695_elements(2)); -- 
    cr_4076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => type_cast_1310_inst_req_1); -- 
    rr_4110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1322_load_0_req_0); -- 
    cr_4057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1306_load_0_req_1); -- 
    rr_3982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => LOAD_padding_1292_load_0_req_0); -- 
    rr_4160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1334_load_0_req_0); -- 
    rr_3949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1289_load_0_req_0); -- 
    cr_4012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => type_cast_1296_inst_req_1); -- 
    cr_3915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => type_cast_1277_inst_req_1); -- 
    rr_3835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1263_load_0_req_0); -- 
    cr_4221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1346_load_0_req_1); -- 
    cr_3846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1263_load_0_req_1); -- 
    rr_4210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1346_load_0_req_0); -- 
    cr_4171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1334_load_0_req_1); -- 
    cr_3960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1289_load_0_req_1); -- 
    rr_4046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1306_load_0_req_0); -- 
    cr_3896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1273_load_0_req_1); -- 
    cr_3993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => LOAD_padding_1292_load_0_req_1); -- 
    cr_4121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1322_load_0_req_1); -- 
    rr_3885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1273_load_0_req_0); -- 
    rr_3785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1251_load_0_req_0); -- 
    cr_3796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1251_load_0_req_1); -- 
    rr_4260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1364_load_0_req_0); -- 
    cr_4271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(2), ack => ptr_deref_1364_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Sample/word_access_start/word_0/ra
      -- 
    ra_3786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1251_load_0_ack_0, ack => convTransposeA_CP_3695_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	29 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Update/ptr_deref_1251_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Update/ptr_deref_1251_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Update/ptr_deref_1251_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1251_Update/ptr_deref_1251_Merge/merge_ack
      -- 
    ca_3797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1251_load_0_ack_1, ack => convTransposeA_CP_3695_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Sample/word_access_start/$exit
      -- 
    ra_3836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1263_load_0_ack_0, ack => convTransposeA_CP_3695_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	29 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Update/ptr_deref_1263_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Update/ptr_deref_1263_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Update/ptr_deref_1263_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Update/ptr_deref_1263_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1263_update_completed_
      -- 
    ca_3847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1263_load_0_ack_1, ack => convTransposeA_CP_3695_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Sample/word_access_start/word_0/$exit
      -- 
    ra_3886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1273_load_0_ack_0, ack => convTransposeA_CP_3695_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Update/ptr_deref_1273_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1277_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Update/ptr_deref_1273_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1277_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1277_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Update/ptr_deref_1273_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Update/ptr_deref_1273_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1273_Update/$exit
      -- 
    ca_3897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1273_load_0_ack_1, ack => convTransposeA_CP_3695_elements(8)); -- 
    rr_3910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(8), ack => type_cast_1277_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1277_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1277_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1277_Sample/$exit
      -- 
    ra_3911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1277_inst_ack_0, ack => convTransposeA_CP_3695_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	29 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1277_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1277_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1277_update_completed_
      -- 
    ca_3916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1277_inst_ack_1, ack => convTransposeA_CP_3695_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Sample/word_access_start/word_0/ra
      -- CP-element group 11: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Sample/word_access_start/word_0/$exit
      -- 
    ra_3950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1289_load_0_ack_0, ack => convTransposeA_CP_3695_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Update/ptr_deref_1289_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Update/ptr_deref_1289_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Update/ptr_deref_1289_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_Update/ptr_deref_1289_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1289_update_completed_
      -- 
    ca_3961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1289_load_0_ack_1, ack => convTransposeA_CP_3695_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Sample/word_access_start/word_0/ra
      -- CP-element group 13: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_sample_completed_
      -- 
    ra_3983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1292_load_0_ack_0, ack => convTransposeA_CP_3695_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (12) 
      -- CP-element group 14: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1296_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1296_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1296_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Update/LOAD_padding_1292_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Update/LOAD_padding_1292_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Update/LOAD_padding_1292_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Update/LOAD_padding_1292_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/LOAD_padding_1292_Update/word_access_complete/$exit
      -- 
    ca_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1292_load_0_ack_1, ack => convTransposeA_CP_3695_elements(14)); -- 
    rr_4007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(14), ack => type_cast_1296_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1296_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1296_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1296_sample_completed_
      -- 
    ra_4008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1296_inst_ack_0, ack => convTransposeA_CP_3695_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1296_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1296_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1296_update_completed_
      -- 
    ca_4013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1296_inst_ack_1, ack => convTransposeA_CP_3695_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Sample/word_access_start/word_0/ra
      -- CP-element group 17: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Sample/word_access_start/$exit
      -- 
    ra_4047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1306_load_0_ack_0, ack => convTransposeA_CP_3695_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (12) 
      -- CP-element group 18: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Update/ptr_deref_1306_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Update/ptr_deref_1306_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Update/ptr_deref_1306_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1310_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Update/ptr_deref_1306_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1306_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1310_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1310_Sample/rr
      -- 
    ca_4058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1306_load_0_ack_1, ack => convTransposeA_CP_3695_elements(18)); -- 
    rr_4071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(18), ack => type_cast_1310_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1310_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1310_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1310_Sample/ra
      -- 
    ra_4072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1310_inst_ack_0, ack => convTransposeA_CP_3695_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	29 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1310_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1310_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/type_cast_1310_Update/ca
      -- 
    ca_4077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1310_inst_ack_1, ack => convTransposeA_CP_3695_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Sample/word_access_start/word_0/ra
      -- CP-element group 21: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Sample/$exit
      -- 
    ra_4111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1322_load_0_ack_0, ack => convTransposeA_CP_3695_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	29 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Update/ptr_deref_1322_Merge/merge_ack
      -- CP-element group 22: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Update/ptr_deref_1322_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Update/ptr_deref_1322_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Update/ptr_deref_1322_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1322_Update/$exit
      -- 
    ca_4122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1322_load_0_ack_1, ack => convTransposeA_CP_3695_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Sample/word_access_start/word_0/ra
      -- CP-element group 23: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_sample_completed_
      -- 
    ra_4161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1334_load_0_ack_0, ack => convTransposeA_CP_3695_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Update/ptr_deref_1334_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Update/ptr_deref_1334_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Update/ptr_deref_1334_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_Update/ptr_deref_1334_Merge/merge_ack
      -- CP-element group 24: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1334_update_completed_
      -- 
    ca_4172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1334_load_0_ack_1, ack => convTransposeA_CP_3695_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Sample/word_access_start/word_0/ra
      -- CP-element group 25: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Sample/word_access_start/$exit
      -- 
    ra_4211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1346_load_0_ack_0, ack => convTransposeA_CP_3695_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Update/ptr_deref_1346_Merge/merge_ack
      -- CP-element group 26: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Update/ptr_deref_1346_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Update/ptr_deref_1346_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1346_Update/ptr_deref_1346_Merge/$exit
      -- 
    ca_4222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1346_load_0_ack_1, ack => convTransposeA_CP_3695_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Sample/word_access_start/word_0/ra
      -- 
    ra_4261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1364_load_0_ack_0, ack => convTransposeA_CP_3695_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Update/ptr_deref_1364_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Update/ptr_deref_1364_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Update/ptr_deref_1364_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/ptr_deref_1364_Update/ptr_deref_1364_Merge/merge_ack
      -- 
    ca_4272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1364_load_0_ack_1, ack => convTransposeA_CP_3695_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  place  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	22 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	26 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	4 
    -- CP-element group 29: 	6 
    -- CP-element group 29: 	10 
    -- CP-element group 29: 	12 
    -- CP-element group 29: 	16 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	69 
    -- CP-element group 29: 	70 
    -- CP-element group 29:  members (8) 
      -- CP-element group 29: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371__exit__
      -- CP-element group 29: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter
      -- CP-element group 29: 	 branch_block_stmt_1236/assign_stmt_1248_to_assign_stmt_1371/$exit
      -- CP-element group 29: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/$entry
      -- CP-element group 29: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/$entry
      -- CP-element group 29: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/$entry
      -- 
    convTransposeA_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeA_CP_3695_elements(20) & convTransposeA_CP_3695_elements(22) & convTransposeA_CP_3695_elements(24) & convTransposeA_CP_3695_elements(26) & convTransposeA_CP_3695_elements(28) & convTransposeA_CP_3695_elements(4) & convTransposeA_CP_3695_elements(6) & convTransposeA_CP_3695_elements(10) & convTransposeA_CP_3695_elements(12) & convTransposeA_CP_3695_elements(16);
      gj_convTransposeA_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3695_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	82 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1393_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1393_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1393_Sample/ra
      -- 
    ra_4289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1393_inst_ack_0, ack => convTransposeA_CP_3695_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	82 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1393_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1393_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1393_Update/ca
      -- 
    ca_4294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1393_inst_ack_1, ack => convTransposeA_CP_3695_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	82 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1398_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1398_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1398_Sample/ra
      -- 
    ra_4303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1398_inst_ack_0, ack => convTransposeA_CP_3695_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	82 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1398_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1398_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1398_Update/ca
      -- 
    ca_4308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1398_inst_ack_1, ack => convTransposeA_CP_3695_elements(33)); -- 
    -- CP-element group 34:  join  transition  place  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	86 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501__exit__
      -- CP-element group 34: 	 branch_block_stmt_1236/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 34: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/$exit
      -- CP-element group 34: 	 branch_block_stmt_1236/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_1236/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1504/$entry
      -- CP-element group 34: 	 branch_block_stmt_1236/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/$entry
      -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3695_elements(31) & convTransposeA_CP_3695_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3695_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	88 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1520_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1520_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1520_Sample/ra
      -- 
    ra_4320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1520_inst_ack_0, ack => convTransposeA_CP_3695_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	88 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	45 
    -- CP-element group 36:  members (9) 
      -- CP-element group 36: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1520_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1520_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1520_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1551_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1551_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1551_Sample/rr
      -- CP-element group 36: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1582_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1582_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1582_Sample/rr
      -- 
    ca_4325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1520_inst_ack_1, ack => convTransposeA_CP_3695_elements(36)); -- 
    rr_4333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(36), ack => type_cast_1551_inst_req_0); -- 
    rr_4443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(36), ack => type_cast_1582_inst_req_0); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1551_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1551_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1551_Sample/ra
      -- 
    ra_4334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1551_inst_ack_0, ack => convTransposeA_CP_3695_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	88 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (16) 
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1551_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1551_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1551_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_index_resized_1
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_index_scaled_1
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_index_computed_1
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_index_resize_1/$entry
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_index_resize_1/$exit
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_index_resize_1/index_resize_req
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_index_resize_1/index_resize_ack
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_index_scale_1/$entry
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_index_scale_1/$exit
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_index_scale_1/scale_rename_req
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_index_scale_1/scale_rename_ack
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_final_index_sum_regn_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_final_index_sum_regn_Sample/req
      -- 
    ca_4339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1551_inst_ack_1, ack => convTransposeA_CP_3695_elements(38)); -- 
    req_4364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(38), ack => array_obj_ref_1557_index_offset_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	56 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_final_index_sum_regn_sample_complete
      -- CP-element group 39: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_final_index_sum_regn_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_final_index_sum_regn_Sample/ack
      -- 
    ack_4365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1557_index_offset_ack_0, ack => convTransposeA_CP_3695_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	88 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (11) 
      -- CP-element group 40: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1558_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_root_address_calculated
      -- CP-element group 40: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_offset_calculated
      -- CP-element group 40: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_final_index_sum_regn_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_final_index_sum_regn_Update/ack
      -- CP-element group 40: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_base_plus_offset/$entry
      -- CP-element group 40: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_base_plus_offset/$exit
      -- CP-element group 40: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_base_plus_offset/sum_rename_req
      -- CP-element group 40: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_base_plus_offset/sum_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1558_request/$entry
      -- CP-element group 40: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1558_request/req
      -- 
    ack_4370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1557_index_offset_ack_1, ack => convTransposeA_CP_3695_elements(40)); -- 
    req_4379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(40), ack => addr_of_1558_final_reg_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1558_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1558_request/$exit
      -- CP-element group 41: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1558_request/ack
      -- 
    ack_4380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1558_final_reg_ack_0, ack => convTransposeA_CP_3695_elements(41)); -- 
    -- CP-element group 42:  join  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	88 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (24) 
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1558_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1558_complete/$exit
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1558_complete/ack
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_base_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_word_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_base_address_resized
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_base_addr_resize/$entry
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_base_addr_resize/$exit
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_base_addr_resize/base_resize_req
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_base_addr_resize/base_resize_ack
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_word_addrgen/$entry
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_word_addrgen/$exit
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_word_addrgen/root_register_req
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_word_addrgen/root_register_ack
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Sample/word_access_start/$entry
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Sample/word_access_start/word_0/$entry
      -- CP-element group 42: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Sample/word_access_start/word_0/rr
      -- 
    ack_4385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1558_final_reg_ack_1, ack => convTransposeA_CP_3695_elements(42)); -- 
    rr_4418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(42), ack => ptr_deref_1562_load_0_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Sample/word_access_start/$exit
      -- CP-element group 43: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Sample/word_access_start/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Sample/word_access_start/word_0/ra
      -- 
    ra_4419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1562_load_0_ack_0, ack => convTransposeA_CP_3695_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	88 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	51 
    -- CP-element group 44:  members (9) 
      -- CP-element group 44: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Update/word_access_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Update/word_access_complete/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Update/word_access_complete/word_0/ca
      -- CP-element group 44: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Update/ptr_deref_1562_Merge/$entry
      -- CP-element group 44: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Update/ptr_deref_1562_Merge/$exit
      -- CP-element group 44: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Update/ptr_deref_1562_Merge/merge_req
      -- CP-element group 44: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Update/ptr_deref_1562_Merge/merge_ack
      -- 
    ca_4430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1562_load_0_ack_1, ack => convTransposeA_CP_3695_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	36 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1582_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1582_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1582_Sample/ra
      -- 
    ra_4444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1582_inst_ack_0, ack => convTransposeA_CP_3695_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	88 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (16) 
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1582_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1582_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1582_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_index_resized_1
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_index_scaled_1
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_index_computed_1
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_index_resize_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_index_resize_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_index_resize_1/index_resize_req
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_index_resize_1/index_resize_ack
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_index_scale_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_index_scale_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_index_scale_1/scale_rename_req
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_index_scale_1/scale_rename_ack
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_final_index_sum_regn_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_final_index_sum_regn_Sample/req
      -- 
    ca_4449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1582_inst_ack_1, ack => convTransposeA_CP_3695_elements(46)); -- 
    req_4474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(46), ack => array_obj_ref_1588_index_offset_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_final_index_sum_regn_sample_complete
      -- CP-element group 47: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_final_index_sum_regn_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_final_index_sum_regn_Sample/ack
      -- 
    ack_4475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1588_index_offset_ack_0, ack => convTransposeA_CP_3695_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	88 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (11) 
      -- CP-element group 48: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1589_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_root_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_offset_calculated
      -- CP-element group 48: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_final_index_sum_regn_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_final_index_sum_regn_Update/ack
      -- CP-element group 48: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_base_plus_offset/$entry
      -- CP-element group 48: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_base_plus_offset/$exit
      -- CP-element group 48: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_base_plus_offset/sum_rename_req
      -- CP-element group 48: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_base_plus_offset/sum_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1589_request/$entry
      -- CP-element group 48: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1589_request/req
      -- 
    ack_4480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1588_index_offset_ack_1, ack => convTransposeA_CP_3695_elements(48)); -- 
    req_4489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(48), ack => addr_of_1589_final_reg_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1589_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1589_request/$exit
      -- CP-element group 49: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1589_request/ack
      -- 
    ack_4490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1589_final_reg_ack_0, ack => convTransposeA_CP_3695_elements(49)); -- 
    -- CP-element group 50:  fork  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	88 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (19) 
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1589_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1589_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1589_complete/ack
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_base_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_word_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_base_address_resized
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_base_addr_resize/$entry
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_base_addr_resize/$exit
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_base_addr_resize/base_resize_req
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_base_addr_resize/base_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_word_addrgen/$entry
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_word_addrgen/$exit
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_word_addrgen/root_register_req
      -- CP-element group 50: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_word_addrgen/root_register_ack
      -- 
    ack_4495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1589_final_reg_ack_1, ack => convTransposeA_CP_3695_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	44 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Sample/ptr_deref_1592_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Sample/ptr_deref_1592_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Sample/ptr_deref_1592_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Sample/ptr_deref_1592_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Sample/word_access_start/word_0/rr
      -- 
    rr_4533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(51), ack => ptr_deref_1592_store_0_req_0); -- 
    convTransposeA_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3695_elements(44) & convTransposeA_CP_3695_elements(50);
      gj_convTransposeA_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3695_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Sample/word_access_start/word_0/ra
      -- 
    ra_4534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1592_store_0_ack_0, ack => convTransposeA_CP_3695_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	88 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Update/word_access_complete/word_0/ca
      -- 
    ca_4545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1592_store_0_ack_1, ack => convTransposeA_CP_3695_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	88 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1598_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1598_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1598_Sample/ra
      -- 
    ra_4554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1598_inst_ack_0, ack => convTransposeA_CP_3695_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	88 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1598_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1598_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1598_Update/ca
      -- 
    ca_4559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1598_inst_ack_1, ack => convTransposeA_CP_3695_elements(55)); -- 
    -- CP-element group 56:  branch  join  transition  place  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: 	47 
    -- CP-element group 56: 	53 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (10) 
      -- CP-element group 56: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610__exit__
      -- CP-element group 56: 	 branch_block_stmt_1236/if_stmt_1611__entry__
      -- CP-element group 56: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/$exit
      -- CP-element group 56: 	 branch_block_stmt_1236/if_stmt_1611_dead_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_1236/if_stmt_1611_eval_test/$entry
      -- CP-element group 56: 	 branch_block_stmt_1236/if_stmt_1611_eval_test/$exit
      -- CP-element group 56: 	 branch_block_stmt_1236/if_stmt_1611_eval_test/branch_req
      -- CP-element group 56: 	 branch_block_stmt_1236/R_cmp_1612_place
      -- CP-element group 56: 	 branch_block_stmt_1236/if_stmt_1611_if_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_1236/if_stmt_1611_else_link/$entry
      -- 
    branch_req_4567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(56), ack => if_stmt_1611_branch_req_0); -- 
    convTransposeA_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3695_elements(39) & convTransposeA_CP_3695_elements(47) & convTransposeA_CP_3695_elements(53) & convTransposeA_CP_3695_elements(55);
      gj_convTransposeA_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3695_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	83 
    -- CP-element group 57: 	84 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_1236/merge_stmt_1617__exit__
      -- CP-element group 57: 	 branch_block_stmt_1236/assign_stmt_1623__entry__
      -- CP-element group 57: 	 branch_block_stmt_1236/assign_stmt_1623__exit__
      -- CP-element group 57: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody
      -- CP-element group 57: 	 branch_block_stmt_1236/if_stmt_1611_if_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_1236/if_stmt_1611_if_link/if_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_1236/whilex_xbody_ifx_xthen
      -- CP-element group 57: 	 branch_block_stmt_1236/assign_stmt_1623/$entry
      -- CP-element group 57: 	 branch_block_stmt_1236/assign_stmt_1623/$exit
      -- CP-element group 57: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/$entry
      -- CP-element group 57: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/$entry
      -- CP-element group 57: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/$entry
      -- CP-element group 57: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/$entry
      -- CP-element group 57: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1236/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1236/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_1236/merge_stmt_1617_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1236/merge_stmt_1617_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_1236/merge_stmt_1617_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_1236/merge_stmt_1617_PhiAck/dummy
      -- 
    if_choice_transition_4572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1611_branch_ack_1, ack => convTransposeA_CP_3695_elements(57)); -- 
    rr_4755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(57), ack => type_cast_1510_inst_req_0); -- 
    cr_4760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(57), ack => type_cast_1510_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	62 
    -- CP-element group 58: 	64 
    -- CP-element group 58:  members (24) 
      -- CP-element group 58: 	 branch_block_stmt_1236/merge_stmt_1625__exit__
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667__entry__
      -- CP-element group 58: 	 branch_block_stmt_1236/if_stmt_1611_else_link/$exit
      -- CP-element group 58: 	 branch_block_stmt_1236/if_stmt_1611_else_link/else_choice_transition
      -- CP-element group 58: 	 branch_block_stmt_1236/whilex_xbody_ifx_xelse
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/$entry
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1635_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1635_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1635_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1635_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1635_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1635_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1644_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1644_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1644_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1661_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1661_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1661_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1236/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1236/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 58: 	 branch_block_stmt_1236/merge_stmt_1625_PhiReqMerge
      -- CP-element group 58: 	 branch_block_stmt_1236/merge_stmt_1625_PhiAck/$entry
      -- CP-element group 58: 	 branch_block_stmt_1236/merge_stmt_1625_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1236/merge_stmt_1625_PhiAck/dummy
      -- 
    else_choice_transition_4576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1611_branch_ack_0, ack => convTransposeA_CP_3695_elements(58)); -- 
    rr_4592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(58), ack => type_cast_1635_inst_req_0); -- 
    cr_4597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(58), ack => type_cast_1635_inst_req_1); -- 
    cr_4611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(58), ack => type_cast_1644_inst_req_1); -- 
    cr_4625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(58), ack => type_cast_1661_inst_req_1); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1635_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1635_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1635_Sample/ra
      -- 
    ra_4593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1635_inst_ack_0, ack => convTransposeA_CP_3695_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1635_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1635_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1635_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1644_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1644_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1644_Sample/rr
      -- 
    ca_4598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1635_inst_ack_1, ack => convTransposeA_CP_3695_elements(60)); -- 
    rr_4606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(60), ack => type_cast_1644_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1644_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1644_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1644_Sample/ra
      -- 
    ra_4607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1644_inst_ack_0, ack => convTransposeA_CP_3695_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	58 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1644_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1644_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1644_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1661_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1661_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1661_Sample/rr
      -- 
    ca_4612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1644_inst_ack_1, ack => convTransposeA_CP_3695_elements(62)); -- 
    rr_4620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(62), ack => type_cast_1661_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1661_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1661_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1661_Sample/ra
      -- 
    ra_4621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1661_inst_ack_0, ack => convTransposeA_CP_3695_elements(63)); -- 
    -- CP-element group 64:  branch  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	58 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (13) 
      -- CP-element group 64: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667__exit__
      -- CP-element group 64: 	 branch_block_stmt_1236/if_stmt_1668__entry__
      -- CP-element group 64: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/$exit
      -- CP-element group 64: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1661_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1661_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1236/assign_stmt_1631_to_assign_stmt_1667/type_cast_1661_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_1236/if_stmt_1668_dead_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_1236/if_stmt_1668_eval_test/$entry
      -- CP-element group 64: 	 branch_block_stmt_1236/if_stmt_1668_eval_test/$exit
      -- CP-element group 64: 	 branch_block_stmt_1236/if_stmt_1668_eval_test/branch_req
      -- CP-element group 64: 	 branch_block_stmt_1236/R_cmp77_1669_place
      -- CP-element group 64: 	 branch_block_stmt_1236/if_stmt_1668_if_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_1236/if_stmt_1668_else_link/$entry
      -- 
    ca_4626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1661_inst_ack_1, ack => convTransposeA_CP_3695_elements(64)); -- 
    branch_req_4634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(64), ack => if_stmt_1668_branch_req_0); -- 
    -- CP-element group 65:  merge  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (15) 
      -- CP-element group 65: 	 branch_block_stmt_1236/merge_stmt_1674__exit__
      -- CP-element group 65: 	 branch_block_stmt_1236/assign_stmt_1678__entry__
      -- CP-element group 65: 	 branch_block_stmt_1236/if_stmt_1668_if_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_1236/if_stmt_1668_if_link/if_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1236/ifx_xelse_whilex_xend
      -- CP-element group 65: 	 branch_block_stmt_1236/assign_stmt_1678/$entry
      -- CP-element group 65: 	 branch_block_stmt_1236/assign_stmt_1678/WPIPE_Block0_done_1676_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_1236/assign_stmt_1678/WPIPE_Block0_done_1676_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1236/assign_stmt_1678/WPIPE_Block0_done_1676_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_1236/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1236/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_1236/merge_stmt_1674_PhiReqMerge
      -- CP-element group 65: 	 branch_block_stmt_1236/merge_stmt_1674_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_1236/merge_stmt_1674_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_1236/merge_stmt_1674_PhiAck/dummy
      -- 
    if_choice_transition_4639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1668_branch_ack_1, ack => convTransposeA_CP_3695_elements(65)); -- 
    req_4656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(65), ack => WPIPE_Block0_done_1676_inst_req_0); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	72 
    -- CP-element group 66: 	73 
    -- CP-element group 66: 	75 
    -- CP-element group 66: 	76 
    -- CP-element group 66:  members (20) 
      -- CP-element group 66: 	 branch_block_stmt_1236/if_stmt_1668_else_link/$exit
      -- CP-element group 66: 	 branch_block_stmt_1236/if_stmt_1668_else_link/else_choice_transition
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/$entry
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/type_cast_1380/$entry
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/type_cast_1380/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/type_cast_1380/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/type_cast_1380/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/type_cast_1380/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/type_cast_1380/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/$entry
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1387/$entry
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1387/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1387/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1387/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1387/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1387/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1668_branch_ack_0, ack => convTransposeA_CP_3695_elements(66)); -- 
    rr_4700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(66), ack => type_cast_1380_inst_req_0); -- 
    cr_4705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(66), ack => type_cast_1380_inst_req_1); -- 
    rr_4723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(66), ack => type_cast_1387_inst_req_0); -- 
    cr_4728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(66), ack => type_cast_1387_inst_req_1); -- 
    -- CP-element group 67:  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_1236/assign_stmt_1678/WPIPE_Block0_done_1676_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1236/assign_stmt_1678/WPIPE_Block0_done_1676_update_start_
      -- CP-element group 67: 	 branch_block_stmt_1236/assign_stmt_1678/WPIPE_Block0_done_1676_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1236/assign_stmt_1678/WPIPE_Block0_done_1676_Sample/ack
      -- CP-element group 67: 	 branch_block_stmt_1236/assign_stmt_1678/WPIPE_Block0_done_1676_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_1236/assign_stmt_1678/WPIPE_Block0_done_1676_Update/req
      -- 
    ack_4657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1676_inst_ack_0, ack => convTransposeA_CP_3695_elements(67)); -- 
    req_4661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(67), ack => WPIPE_Block0_done_1676_inst_req_1); -- 
    -- CP-element group 68:  transition  place  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 $exit
      -- CP-element group 68: 	 branch_block_stmt_1236/$exit
      -- CP-element group 68: 	 branch_block_stmt_1236/branch_block_stmt_1236__exit__
      -- CP-element group 68: 	 branch_block_stmt_1236/assign_stmt_1678__exit__
      -- CP-element group 68: 	 branch_block_stmt_1236/return__
      -- CP-element group 68: 	 branch_block_stmt_1236/merge_stmt_1680__exit__
      -- CP-element group 68: 	 branch_block_stmt_1236/assign_stmt_1678/$exit
      -- CP-element group 68: 	 branch_block_stmt_1236/assign_stmt_1678/WPIPE_Block0_done_1676_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_1236/assign_stmt_1678/WPIPE_Block0_done_1676_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1236/assign_stmt_1678/WPIPE_Block0_done_1676_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_1236/return___PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_1236/return___PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_1236/merge_stmt_1680_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_1236/merge_stmt_1680_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_1236/merge_stmt_1680_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_1236/merge_stmt_1680_PhiAck/dummy
      -- 
    ack_4662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1676_inst_ack_1, ack => convTransposeA_CP_3695_elements(68)); -- 
    -- CP-element group 69:  transition  output  delay-element  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	29 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/$exit
      -- CP-element group 69: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/type_cast_1378_konst_delay_trans
      -- CP-element group 69: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_req
      -- 
    phi_stmt_1374_req_4673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1374_req_4673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(69), ack => phi_stmt_1374_req_0); -- 
    -- Element group convTransposeA_CP_3695_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => convTransposeA_CP_3695_elements(29), ack => convTransposeA_CP_3695_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  transition  output  delay-element  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	29 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/$exit
      -- CP-element group 70: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1385_konst_delay_trans
      -- CP-element group 70: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_req
      -- 
    phi_stmt_1381_req_4681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1381_req_4681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(70), ack => phi_stmt_1381_req_0); -- 
    -- Element group convTransposeA_CP_3695_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => convTransposeA_CP_3695_elements(29), ack => convTransposeA_CP_3695_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  transition  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	79 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1236/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3695_elements(69) & convTransposeA_CP_3695_elements(70);
      gj_convTransposeA_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3695_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	66 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/type_cast_1380/SplitProtocol/Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/type_cast_1380/SplitProtocol/Sample/ra
      -- 
    ra_4701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1380_inst_ack_0, ack => convTransposeA_CP_3695_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	66 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/type_cast_1380/SplitProtocol/Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/type_cast_1380/SplitProtocol/Update/ca
      -- 
    ca_4706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1380_inst_ack_1, ack => convTransposeA_CP_3695_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	78 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/$exit
      -- CP-element group 74: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/type_cast_1380/$exit
      -- CP-element group 74: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_sources/type_cast_1380/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1374/phi_stmt_1374_req
      -- 
    phi_stmt_1374_req_4707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1374_req_4707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(74), ack => phi_stmt_1374_req_1); -- 
    convTransposeA_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3695_elements(72) & convTransposeA_CP_3695_elements(73);
      gj_convTransposeA_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3695_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	66 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1387/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1387/SplitProtocol/Sample/ra
      -- 
    ra_4724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1387_inst_ack_0, ack => convTransposeA_CP_3695_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	66 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1387/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1387/SplitProtocol/Update/ca
      -- 
    ca_4729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1387_inst_ack_1, ack => convTransposeA_CP_3695_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/$exit
      -- CP-element group 77: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1387/$exit
      -- CP-element group 77: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1387/SplitProtocol/$exit
      -- CP-element group 77: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1381/phi_stmt_1381_req
      -- 
    phi_stmt_1381_req_4730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1381_req_4730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(77), ack => phi_stmt_1381_req_1); -- 
    convTransposeA_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3695_elements(75) & convTransposeA_CP_3695_elements(76);
      gj_convTransposeA_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3695_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	74 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1236/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3695_elements(74) & convTransposeA_CP_3695_elements(77);
      gj_convTransposeA_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3695_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  merge  fork  transition  place  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	71 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1236/merge_stmt_1373_PhiReqMerge
      -- CP-element group 79: 	 branch_block_stmt_1236/merge_stmt_1373_PhiAck/$entry
      -- 
    convTransposeA_CP_3695_elements(79) <= OrReduce(convTransposeA_CP_3695_elements(71) & convTransposeA_CP_3695_elements(78));
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1236/merge_stmt_1373_PhiAck/phi_stmt_1374_ack
      -- 
    phi_stmt_1374_ack_4735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1374_ack_0, ack => convTransposeA_CP_3695_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1236/merge_stmt_1373_PhiAck/phi_stmt_1381_ack
      -- 
    phi_stmt_1381_ack_4736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1381_ack_0, ack => convTransposeA_CP_3695_elements(81)); -- 
    -- CP-element group 82:  join  fork  transition  place  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	30 
    -- CP-element group 82: 	31 
    -- CP-element group 82: 	32 
    -- CP-element group 82: 	33 
    -- CP-element group 82:  members (16) 
      -- CP-element group 82: 	 branch_block_stmt_1236/merge_stmt_1373__exit__
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501__entry__
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/$entry
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1393_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1393_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1393_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1393_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1393_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1393_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1398_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1398_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1398_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1398_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1398_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1236/assign_stmt_1394_to_assign_stmt_1501/type_cast_1398_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1236/merge_stmt_1373_PhiAck/$exit
      -- 
    rr_4288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(82), ack => type_cast_1393_inst_req_0); -- 
    cr_4293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(82), ack => type_cast_1393_inst_req_1); -- 
    rr_4302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(82), ack => type_cast_1398_inst_req_0); -- 
    cr_4307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(82), ack => type_cast_1398_inst_req_1); -- 
    convTransposeA_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3695_elements(80) & convTransposeA_CP_3695_elements(81);
      gj_convTransposeA_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3695_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	57 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Sample/ra
      -- 
    ra_4756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1510_inst_ack_0, ack => convTransposeA_CP_3695_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	57 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Update/ca
      -- 
    ca_4761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1510_inst_ack_1, ack => convTransposeA_CP_3695_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/$exit
      -- CP-element group 85: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/$exit
      -- CP-element group 85: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/$exit
      -- CP-element group 85: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/$exit
      -- CP-element group 85: 	 branch_block_stmt_1236/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_req
      -- 
    phi_stmt_1504_req_4762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1504_req_4762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(85), ack => phi_stmt_1504_req_1); -- 
    convTransposeA_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3695_elements(83) & convTransposeA_CP_3695_elements(84);
      gj_convTransposeA_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3695_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  output  delay-element  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	34 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1236/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_1236/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1504/$exit
      -- CP-element group 86: 	 branch_block_stmt_1236/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1236/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1508_konst_delay_trans
      -- CP-element group 86: 	 branch_block_stmt_1236/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1504/phi_stmt_1504_req
      -- 
    phi_stmt_1504_req_4773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1504_req_4773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(86), ack => phi_stmt_1504_req_0); -- 
    -- Element group convTransposeA_CP_3695_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => convTransposeA_CP_3695_elements(34), ack => convTransposeA_CP_3695_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  merge  transition  place  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1236/merge_stmt_1503_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_1236/merge_stmt_1503_PhiAck/$entry
      -- 
    convTransposeA_CP_3695_elements(87) <= OrReduce(convTransposeA_CP_3695_elements(85) & convTransposeA_CP_3695_elements(86));
    -- CP-element group 88:  fork  transition  place  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	35 
    -- CP-element group 88: 	36 
    -- CP-element group 88: 	38 
    -- CP-element group 88: 	40 
    -- CP-element group 88: 	42 
    -- CP-element group 88: 	44 
    -- CP-element group 88: 	46 
    -- CP-element group 88: 	48 
    -- CP-element group 88: 	50 
    -- CP-element group 88: 	53 
    -- CP-element group 88: 	54 
    -- CP-element group 88: 	55 
    -- CP-element group 88:  members (45) 
      -- CP-element group 88: 	 branch_block_stmt_1236/merge_stmt_1503__exit__
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610__entry__
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1520_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1520_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1520_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1520_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1520_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1520_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1551_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1551_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1551_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1558_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_final_index_sum_regn_update_start
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_final_index_sum_regn_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1557_final_index_sum_regn_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1558_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1558_complete/req
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1562_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1582_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1582_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1582_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1589_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_final_index_sum_regn_update_start
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_final_index_sum_regn_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/array_obj_ref_1588_final_index_sum_regn_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1589_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/addr_of_1589_complete/req
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/ptr_deref_1592_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1598_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1598_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1598_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1598_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1598_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1236/assign_stmt_1517_to_assign_stmt_1610/type_cast_1598_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1236/merge_stmt_1503_PhiAck/$exit
      -- CP-element group 88: 	 branch_block_stmt_1236/merge_stmt_1503_PhiAck/phi_stmt_1504_ack
      -- 
    phi_stmt_1504_ack_4778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1504_ack_0, ack => convTransposeA_CP_3695_elements(88)); -- 
    rr_4319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(88), ack => type_cast_1520_inst_req_0); -- 
    cr_4324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(88), ack => type_cast_1520_inst_req_1); -- 
    cr_4338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(88), ack => type_cast_1551_inst_req_1); -- 
    req_4369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(88), ack => array_obj_ref_1557_index_offset_req_1); -- 
    req_4384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(88), ack => addr_of_1558_final_reg_req_1); -- 
    cr_4429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(88), ack => ptr_deref_1562_load_0_req_1); -- 
    cr_4448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(88), ack => type_cast_1582_inst_req_1); -- 
    req_4479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(88), ack => array_obj_ref_1588_index_offset_req_1); -- 
    req_4494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(88), ack => addr_of_1589_final_reg_req_1); -- 
    cr_4544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(88), ack => ptr_deref_1592_store_0_req_1); -- 
    rr_4553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(88), ack => type_cast_1598_inst_req_0); -- 
    cr_4558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3695_elements(88), ack => type_cast_1598_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1463_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1484_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1544_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1576_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_1292_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_1292_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom52_1587_resized : std_logic_vector(13 downto 0);
    signal R_idxprom52_1587_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1556_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1556_scaled : std_logic_vector(13 downto 0);
    signal add16_1424 : std_logic_vector(31 downto 0);
    signal add27_1439 : std_logic_vector(31 downto 0);
    signal add42_1496 : std_logic_vector(31 downto 0);
    signal add44_1531 : std_logic_vector(31 downto 0);
    signal add57_1605 : std_logic_vector(31 downto 0);
    signal add8_1526 : std_logic_vector(31 downto 0);
    signal add_1409 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1557_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1557_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1557_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1557_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1557_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1557_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1588_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1588_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1588_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1588_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1588_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1588_root_address : std_logic_vector(13 downto 0);
    signal arrayidx53_1590 : std_logic_vector(31 downto 0);
    signal arrayidx_1559 : std_logic_vector(31 downto 0);
    signal call_1239 : std_logic_vector(15 downto 0);
    signal cmp68_1641 : std_logic_vector(0 downto 0);
    signal cmp77_1667 : std_logic_vector(0 downto 0);
    signal cmp_1610 : std_logic_vector(0 downto 0);
    signal conv13_1278 : std_logic_vector(31 downto 0);
    signal conv18_1297 : std_logic_vector(31 downto 0);
    signal conv24_1311 : std_logic_vector(31 downto 0);
    signal conv37_1465 : std_logic_vector(31 downto 0);
    signal conv3_1394 : std_logic_vector(31 downto 0);
    signal conv40_1486 : std_logic_vector(31 downto 0);
    signal conv56_1599 : std_logic_vector(31 downto 0);
    signal conv66_1636 : std_logic_vector(31 downto 0);
    signal conv6_1399 : std_logic_vector(31 downto 0);
    signal conv74_1662 : std_logic_vector(31 downto 0);
    signal conv90_1521 : std_logic_vector(31 downto 0);
    signal div76_1371 : std_logic_vector(31 downto 0);
    signal div_1353 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1361 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1248 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1260 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1270 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1286 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1303 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1319 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1331 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1343 : std_logic_vector(31 downto 0);
    signal idxprom52_1583 : std_logic_vector(63 downto 0);
    signal idxprom_1552 : std_logic_vector(63 downto 0);
    signal inc72_1645 : std_logic_vector(15 downto 0);
    signal inc72x_xinput_dim0x_x2_1650 : std_logic_vector(15 downto 0);
    signal inc_1631 : std_logic_vector(15 downto 0);
    signal indvar_1504 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1623 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1381 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1374 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1657 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1517 : std_logic_vector(15 downto 0);
    signal mul14_1419 : std_logic_vector(31 downto 0);
    signal mul25_1434 : std_logic_vector(31 downto 0);
    signal mul41_1491 : std_logic_vector(31 downto 0);
    signal mul43_1501 : std_logic_vector(31 downto 0);
    signal mul7_1414 : std_logic_vector(31 downto 0);
    signal mul_1404 : std_logic_vector(31 downto 0);
    signal ptr_deref_1251_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1251_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1251_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1251_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1251_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1263_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1263_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1263_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1263_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1263_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1273_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1273_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1273_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1273_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1273_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1289_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1289_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1289_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1289_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1289_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1306_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1306_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1306_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1306_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1306_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1322_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1322_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1322_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1322_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1322_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1334_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1334_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1334_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1334_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1334_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1346_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1346_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1346_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1346_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1346_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1364_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1364_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1364_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1364_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1364_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1562_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1562_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1562_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1562_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1562_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1592_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1592_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1592_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1592_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1592_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1592_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext91_1477 : std_logic_vector(31 downto 0);
    signal sext93_1537 : std_logic_vector(31 downto 0);
    signal sext94_1569 : std_logic_vector(31 downto 0);
    signal sext_1456 : std_logic_vector(31 downto 0);
    signal shr51_1578 : std_logic_vector(31 downto 0);
    signal shr_1546 : std_logic_vector(31 downto 0);
    signal sub19_1471 : std_logic_vector(31 downto 0);
    signal sub30_1444 : std_logic_vector(31 downto 0);
    signal sub31_1450 : std_logic_vector(31 downto 0);
    signal sub_1429 : std_logic_vector(31 downto 0);
    signal tmp12_1274 : std_logic_vector(15 downto 0);
    signal tmp15_1290 : std_logic_vector(31 downto 0);
    signal tmp17_1293 : std_logic_vector(15 downto 0);
    signal tmp1_1252 : std_logic_vector(31 downto 0);
    signal tmp23_1307 : std_logic_vector(15 downto 0);
    signal tmp26_1323 : std_logic_vector(31 downto 0);
    signal tmp35_1335 : std_logic_vector(31 downto 0);
    signal tmp38_1347 : std_logic_vector(31 downto 0);
    signal tmp48_1563 : std_logic_vector(63 downto 0);
    signal tmp4_1264 : std_logic_vector(31 downto 0);
    signal tmp75_1365 : std_logic_vector(31 downto 0);
    signal type_cast_1351_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1369_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1378_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1380_wire : std_logic_vector(15 downto 0);
    signal type_cast_1385_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1387_wire : std_logic_vector(15 downto 0);
    signal type_cast_1392_wire : std_logic_vector(31 downto 0);
    signal type_cast_1397_wire : std_logic_vector(31 downto 0);
    signal type_cast_1448_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1454_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1459_wire : std_logic_vector(31 downto 0);
    signal type_cast_1462_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1469_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1475_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1480_wire : std_logic_vector(31 downto 0);
    signal type_cast_1483_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1508_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1510_wire : std_logic_vector(15 downto 0);
    signal type_cast_1515_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1535_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1540_wire : std_logic_vector(31 downto 0);
    signal type_cast_1543_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1550_wire : std_logic_vector(63 downto 0);
    signal type_cast_1567_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1572_wire : std_logic_vector(31 downto 0);
    signal type_cast_1575_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1581_wire : std_logic_vector(63 downto 0);
    signal type_cast_1597_wire : std_logic_vector(31 downto 0);
    signal type_cast_1603_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1621_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1629_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1634_wire : std_logic_vector(31 downto 0);
    signal type_cast_1654_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1660_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_1292_word_address_0 <= "0";
    array_obj_ref_1557_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1557_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1557_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1557_resized_base_address <= "00000000000000";
    array_obj_ref_1588_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1588_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1588_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1588_resized_base_address <= "00000000000000";
    iNsTr_10_1361 <= "00000000000000000000000000000010";
    iNsTr_2_1248 <= "00000000000000000000000000000100";
    iNsTr_3_1260 <= "00000000000000000000000000000011";
    iNsTr_4_1270 <= "00000000000000000000000000000000";
    iNsTr_5_1286 <= "00000000000000000000000000000011";
    iNsTr_6_1303 <= "00000000000000000000000000000001";
    iNsTr_7_1319 <= "00000000000000000000000000000100";
    iNsTr_8_1331 <= "00000000000000000000000000000100";
    iNsTr_9_1343 <= "00000000000000000000000000000011";
    ptr_deref_1251_word_offset_0 <= "0000000";
    ptr_deref_1263_word_offset_0 <= "0000000";
    ptr_deref_1273_word_offset_0 <= "0";
    ptr_deref_1289_word_offset_0 <= "0000000";
    ptr_deref_1306_word_offset_0 <= "0";
    ptr_deref_1322_word_offset_0 <= "0000000";
    ptr_deref_1334_word_offset_0 <= "0000000";
    ptr_deref_1346_word_offset_0 <= "0000000";
    ptr_deref_1364_word_offset_0 <= "0000000";
    ptr_deref_1562_word_offset_0 <= "00000000000000";
    ptr_deref_1592_word_offset_0 <= "00000000000000";
    type_cast_1351_wire_constant <= "00000000000000000000000000000001";
    type_cast_1369_wire_constant <= "00000000000000000000000000000001";
    type_cast_1378_wire_constant <= "0000000000000000";
    type_cast_1385_wire_constant <= "0000000000000000";
    type_cast_1448_wire_constant <= "00000000000000000000000000010000";
    type_cast_1454_wire_constant <= "11111111111111110000000000000000";
    type_cast_1462_wire_constant <= "00000000000000000000000000010000";
    type_cast_1469_wire_constant <= "00000000000000000000000000010000";
    type_cast_1475_wire_constant <= "11111111111111110000000000000000";
    type_cast_1483_wire_constant <= "00000000000000000000000000010000";
    type_cast_1508_wire_constant <= "0000000000000000";
    type_cast_1515_wire_constant <= "0000000000000100";
    type_cast_1535_wire_constant <= "00000000000000000000000000010000";
    type_cast_1543_wire_constant <= "00000000000000000000000000010010";
    type_cast_1567_wire_constant <= "00000000000000000000000000010000";
    type_cast_1575_wire_constant <= "00000000000000000000000000010010";
    type_cast_1603_wire_constant <= "00000000000000000000000000000100";
    type_cast_1621_wire_constant <= "0000000000000001";
    type_cast_1629_wire_constant <= "0000000000000001";
    type_cast_1654_wire_constant <= "0000000000000000";
    phi_stmt_1374: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1378_wire_constant & type_cast_1380_wire;
      req <= phi_stmt_1374_req_0 & phi_stmt_1374_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1374",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1374_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1374,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1374
    phi_stmt_1381: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1385_wire_constant & type_cast_1387_wire;
      req <= phi_stmt_1381_req_0 & phi_stmt_1381_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1381",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1381_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1381,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1381
    phi_stmt_1504: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1508_wire_constant & type_cast_1510_wire;
      req <= phi_stmt_1504_req_0 & phi_stmt_1504_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1504",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1504_ack_0,
          idata => idata,
          odata => indvar_1504,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1504
    -- flow-through select operator MUX_1656_inst
    input_dim1x_x2_1657 <= type_cast_1654_wire_constant when (cmp68_1641(0) /=  '0') else inc_1631;
    addr_of_1558_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1558_final_reg_req_0;
      addr_of_1558_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1558_final_reg_req_1;
      addr_of_1558_final_reg_ack_1<= rack(0);
      addr_of_1558_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1558_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1557_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1559,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1589_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1589_final_reg_req_0;
      addr_of_1589_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1589_final_reg_req_1;
      addr_of_1589_final_reg_ack_1<= rack(0);
      addr_of_1589_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1589_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1588_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx53_1590,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1277_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1277_inst_req_0;
      type_cast_1277_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1277_inst_req_1;
      type_cast_1277_inst_ack_1<= rack(0);
      type_cast_1277_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1277_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_1274,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13_1278,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1296_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1296_inst_req_0;
      type_cast_1296_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1296_inst_req_1;
      type_cast_1296_inst_ack_1<= rack(0);
      type_cast_1296_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1296_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp17_1293,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_1297,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1310_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1310_inst_req_0;
      type_cast_1310_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1310_inst_req_1;
      type_cast_1310_inst_ack_1<= rack(0);
      type_cast_1310_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1310_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp23_1307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_1311,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1380_inst_req_0;
      type_cast_1380_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1380_inst_req_1;
      type_cast_1380_inst_ack_1<= rack(0);
      type_cast_1380_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1380_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1657,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1380_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1387_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1387_inst_req_0;
      type_cast_1387_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1387_inst_req_1;
      type_cast_1387_inst_ack_1<= rack(0);
      type_cast_1387_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1387_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc72x_xinput_dim0x_x2_1650,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1387_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1393_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1393_inst_req_0;
      type_cast_1393_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1393_inst_req_1;
      type_cast_1393_inst_ack_1<= rack(0);
      type_cast_1393_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1393_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1392_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_1394,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1398_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1398_inst_req_0;
      type_cast_1398_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1398_inst_req_1;
      type_cast_1398_inst_ack_1<= rack(0);
      type_cast_1398_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1398_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1397_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv6_1399,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1459_inst
    process(sext_1456) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_1456(31 downto 0);
      type_cast_1459_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1464_inst
    process(ASHR_i32_i32_1463_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1463_wire(31 downto 0);
      conv37_1465 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1480_inst
    process(sext91_1477) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext91_1477(31 downto 0);
      type_cast_1480_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1485_inst
    process(ASHR_i32_i32_1484_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1484_wire(31 downto 0);
      conv40_1486 <= tmp_var; -- 
    end process;
    type_cast_1510_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1510_inst_req_0;
      type_cast_1510_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1510_inst_req_1;
      type_cast_1510_inst_ack_1<= rack(0);
      type_cast_1510_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1510_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1623,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1510_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1520_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1520_inst_req_0;
      type_cast_1520_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1520_inst_req_1;
      type_cast_1520_inst_ack_1<= rack(0);
      type_cast_1520_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1520_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1517,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1521,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1540_inst
    process(sext93_1537) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext93_1537(31 downto 0);
      type_cast_1540_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1545_inst
    process(ASHR_i32_i32_1544_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1544_wire(31 downto 0);
      shr_1546 <= tmp_var; -- 
    end process;
    type_cast_1551_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1551_inst_req_0;
      type_cast_1551_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1551_inst_req_1;
      type_cast_1551_inst_ack_1<= rack(0);
      type_cast_1551_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1551_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1550_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1552,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1572_inst
    process(sext94_1569) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext94_1569(31 downto 0);
      type_cast_1572_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1577_inst
    process(ASHR_i32_i32_1576_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1576_wire(31 downto 0);
      shr51_1578 <= tmp_var; -- 
    end process;
    type_cast_1582_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1582_inst_req_0;
      type_cast_1582_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1582_inst_req_1;
      type_cast_1582_inst_ack_1<= rack(0);
      type_cast_1582_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1582_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1581_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom52_1583,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1598_inst_req_0;
      type_cast_1598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1598_inst_req_1;
      type_cast_1598_inst_ack_1<= rack(0);
      type_cast_1598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1598_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1597_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_1599,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1635_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1635_inst_req_0;
      type_cast_1635_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1635_inst_req_1;
      type_cast_1635_inst_ack_1<= rack(0);
      type_cast_1635_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1635_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1634_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1636,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1644_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1644_inst_req_0;
      type_cast_1644_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1644_inst_req_1;
      type_cast_1644_inst_ack_1<= rack(0);
      type_cast_1644_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1644_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp68_1641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc72_1645,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1661_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1661_inst_req_0;
      type_cast_1661_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1661_inst_req_1;
      type_cast_1661_inst_ack_1<= rack(0);
      type_cast_1661_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1661_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1660_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_1662,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1292_gather_scatter
    process(LOAD_padding_1292_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1292_data_0;
      ov(15 downto 0) := iv;
      tmp17_1293 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1557_index_1_rename
    process(R_idxprom_1556_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1556_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1556_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1557_index_1_resize
    process(idxprom_1552) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1552;
      ov := iv(13 downto 0);
      R_idxprom_1556_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1557_root_address_inst
    process(array_obj_ref_1557_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1557_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1557_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1588_index_1_rename
    process(R_idxprom52_1587_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom52_1587_resized;
      ov(13 downto 0) := iv;
      R_idxprom52_1587_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1588_index_1_resize
    process(idxprom52_1583) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom52_1583;
      ov := iv(13 downto 0);
      R_idxprom52_1587_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1588_root_address_inst
    process(array_obj_ref_1588_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1588_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1588_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1251_addr_0
    process(ptr_deref_1251_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1251_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1251_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1251_base_resize
    process(iNsTr_2_1248) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1248;
      ov := iv(6 downto 0);
      ptr_deref_1251_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1251_gather_scatter
    process(ptr_deref_1251_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1251_data_0;
      ov(31 downto 0) := iv;
      tmp1_1252 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1251_root_address_inst
    process(ptr_deref_1251_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1251_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1251_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1263_addr_0
    process(ptr_deref_1263_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1263_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1263_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1263_base_resize
    process(iNsTr_3_1260) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1260;
      ov := iv(6 downto 0);
      ptr_deref_1263_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1263_gather_scatter
    process(ptr_deref_1263_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1263_data_0;
      ov(31 downto 0) := iv;
      tmp4_1264 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1263_root_address_inst
    process(ptr_deref_1263_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1263_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1263_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1273_addr_0
    process(ptr_deref_1273_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1273_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1273_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1273_base_resize
    process(iNsTr_4_1270) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1270;
      ov := iv(0 downto 0);
      ptr_deref_1273_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1273_gather_scatter
    process(ptr_deref_1273_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1273_data_0;
      ov(15 downto 0) := iv;
      tmp12_1274 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1273_root_address_inst
    process(ptr_deref_1273_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1273_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1273_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1289_addr_0
    process(ptr_deref_1289_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1289_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1289_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1289_base_resize
    process(iNsTr_5_1286) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1286;
      ov := iv(6 downto 0);
      ptr_deref_1289_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1289_gather_scatter
    process(ptr_deref_1289_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1289_data_0;
      ov(31 downto 0) := iv;
      tmp15_1290 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1289_root_address_inst
    process(ptr_deref_1289_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1289_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1289_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1306_addr_0
    process(ptr_deref_1306_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1306_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1306_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1306_base_resize
    process(iNsTr_6_1303) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1303;
      ov := iv(0 downto 0);
      ptr_deref_1306_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1306_gather_scatter
    process(ptr_deref_1306_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1306_data_0;
      ov(15 downto 0) := iv;
      tmp23_1307 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1306_root_address_inst
    process(ptr_deref_1306_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1306_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1306_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1322_addr_0
    process(ptr_deref_1322_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1322_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1322_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1322_base_resize
    process(iNsTr_7_1319) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1319;
      ov := iv(6 downto 0);
      ptr_deref_1322_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1322_gather_scatter
    process(ptr_deref_1322_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1322_data_0;
      ov(31 downto 0) := iv;
      tmp26_1323 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1322_root_address_inst
    process(ptr_deref_1322_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1322_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1322_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1334_addr_0
    process(ptr_deref_1334_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1334_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1334_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1334_base_resize
    process(iNsTr_8_1331) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1331;
      ov := iv(6 downto 0);
      ptr_deref_1334_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1334_gather_scatter
    process(ptr_deref_1334_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1334_data_0;
      ov(31 downto 0) := iv;
      tmp35_1335 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1334_root_address_inst
    process(ptr_deref_1334_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1334_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1334_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1346_addr_0
    process(ptr_deref_1346_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1346_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1346_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1346_base_resize
    process(iNsTr_9_1343) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1343;
      ov := iv(6 downto 0);
      ptr_deref_1346_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1346_gather_scatter
    process(ptr_deref_1346_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1346_data_0;
      ov(31 downto 0) := iv;
      tmp38_1347 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1346_root_address_inst
    process(ptr_deref_1346_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1346_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1346_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1364_addr_0
    process(ptr_deref_1364_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1364_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1364_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1364_base_resize
    process(iNsTr_10_1361) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1361;
      ov := iv(6 downto 0);
      ptr_deref_1364_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1364_gather_scatter
    process(ptr_deref_1364_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1364_data_0;
      ov(31 downto 0) := iv;
      tmp75_1365 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1364_root_address_inst
    process(ptr_deref_1364_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1364_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1364_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1562_addr_0
    process(ptr_deref_1562_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1562_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1562_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1562_base_resize
    process(arrayidx_1559) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1559;
      ov := iv(13 downto 0);
      ptr_deref_1562_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1562_gather_scatter
    process(ptr_deref_1562_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1562_data_0;
      ov(63 downto 0) := iv;
      tmp48_1563 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1562_root_address_inst
    process(ptr_deref_1562_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1562_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1562_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1592_addr_0
    process(ptr_deref_1592_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1592_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1592_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1592_base_resize
    process(arrayidx53_1590) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx53_1590;
      ov := iv(13 downto 0);
      ptr_deref_1592_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1592_gather_scatter
    process(tmp48_1563) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp48_1563;
      ov(63 downto 0) := iv;
      ptr_deref_1592_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1592_root_address_inst
    process(ptr_deref_1592_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1592_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1592_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1611_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1610;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1611_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1611_branch_req_0,
          ack0 => if_stmt_1611_branch_ack_0,
          ack1 => if_stmt_1611_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1668_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_1667;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1668_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1668_branch_req_0,
          ack0 => if_stmt_1668_branch_ack_0,
          ack1 => if_stmt_1668_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1622_inst
    process(indvar_1504) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1504, type_cast_1621_wire_constant, tmp_var);
      indvarx_xnext_1623 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1630_inst
    process(input_dim1x_x1x_xph_1374) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1374, type_cast_1629_wire_constant, tmp_var);
      inc_1631 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1649_inst
    process(inc72_1645, input_dim0x_x2x_xph_1381) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc72_1645, input_dim0x_x2x_xph_1381, tmp_var);
      inc72x_xinput_dim0x_x2_1650 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1408_inst
    process(mul_1404, conv3_1394) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_1404, conv3_1394, tmp_var);
      add_1409 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1423_inst
    process(mul14_1419, tmp15_1290) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul14_1419, tmp15_1290, tmp_var);
      add16_1424 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1438_inst
    process(mul25_1434, tmp26_1323) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul25_1434, tmp26_1323, tmp_var);
      add27_1439 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1455_inst
    process(sub31_1450) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub31_1450, type_cast_1454_wire_constant, tmp_var);
      sext_1456 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1476_inst
    process(sub19_1471) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub19_1471, type_cast_1475_wire_constant, tmp_var);
      sext91_1477 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1495_inst
    process(conv37_1465, mul41_1491) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv37_1465, mul41_1491, tmp_var);
      add42_1496 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1525_inst
    process(mul7_1414, conv90_1521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul7_1414, conv90_1521, tmp_var);
      add8_1526 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1530_inst
    process(mul43_1501, conv90_1521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul43_1501, conv90_1521, tmp_var);
      add44_1531 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1604_inst
    process(conv56_1599) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv56_1599, type_cast_1603_wire_constant, tmp_var);
      add57_1605 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1463_inst
    process(type_cast_1459_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1459_wire, type_cast_1462_wire_constant, tmp_var);
      ASHR_i32_i32_1463_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1484_inst
    process(type_cast_1480_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1480_wire, type_cast_1483_wire_constant, tmp_var);
      ASHR_i32_i32_1484_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1544_inst
    process(type_cast_1540_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1540_wire, type_cast_1543_wire_constant, tmp_var);
      ASHR_i32_i32_1544_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1576_inst
    process(type_cast_1572_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1572_wire, type_cast_1575_wire_constant, tmp_var);
      ASHR_i32_i32_1576_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1640_inst
    process(conv66_1636, div_1353) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv66_1636, div_1353, tmp_var);
      cmp68_1641 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1666_inst
    process(conv74_1662, div76_1371) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv74_1662, div76_1371, tmp_var);
      cmp77_1667 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1352_inst
    process(tmp4_1264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1264, type_cast_1351_wire_constant, tmp_var);
      div_1353 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1370_inst
    process(tmp75_1365) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp75_1365, type_cast_1369_wire_constant, tmp_var);
      div76_1371 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1516_inst
    process(indvar_1504) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1504, type_cast_1515_wire_constant, tmp_var);
      input_dim2x_x1_1517 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1403_inst
    process(tmp4_1264, conv6_1399) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp4_1264, conv6_1399, tmp_var);
      mul_1404 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1413_inst
    process(add_1409, tmp1_1252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1409, tmp1_1252, tmp_var);
      mul7_1414 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1418_inst
    process(conv13_1278, conv6_1399) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv13_1278, conv6_1399, tmp_var);
      mul14_1419 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1433_inst
    process(conv24_1311, conv3_1394) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv24_1311, conv3_1394, tmp_var);
      mul25_1434 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1490_inst
    process(tmp38_1347, conv40_1486) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp38_1347, conv40_1486, tmp_var);
      mul41_1491 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1500_inst
    process(add42_1496, tmp35_1335) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add42_1496, tmp35_1335, tmp_var);
      mul43_1501 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1449_inst
    process(sub30_1444) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub30_1444, type_cast_1448_wire_constant, tmp_var);
      sub31_1450 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1470_inst
    process(sub_1429) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_1429, type_cast_1469_wire_constant, tmp_var);
      sub19_1471 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1536_inst
    process(add8_1526) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add8_1526, type_cast_1535_wire_constant, tmp_var);
      sext93_1537 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1568_inst
    process(add44_1531) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add44_1531, type_cast_1567_wire_constant, tmp_var);
      sext94_1569 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1428_inst
    process(add16_1424, conv18_1297) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add16_1424, conv18_1297, tmp_var);
      sub_1429 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1443_inst
    process(add27_1439, conv18_1297) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add27_1439, conv18_1297, tmp_var);
      sub30_1444 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1609_inst
    process(add57_1605, tmp1_1252) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add57_1605, tmp1_1252, tmp_var);
      cmp_1610 <= tmp_var; --
    end process;
    -- shared split operator group (34) : array_obj_ref_1557_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1556_scaled;
      array_obj_ref_1557_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1557_index_offset_req_0;
      array_obj_ref_1557_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1557_index_offset_req_1;
      array_obj_ref_1557_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_1588_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom52_1587_scaled;
      array_obj_ref_1588_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1588_index_offset_req_0;
      array_obj_ref_1588_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1588_index_offset_req_1;
      array_obj_ref_1588_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- unary operator type_cast_1392_inst
    process(input_dim1x_x1x_xph_1374) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_1374, tmp_var);
      type_cast_1392_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1397_inst
    process(input_dim0x_x2x_xph_1381) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_1381, tmp_var);
      type_cast_1397_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1550_inst
    process(shr_1546) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1546, tmp_var);
      type_cast_1550_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1581_inst
    process(shr51_1578) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr51_1578, tmp_var);
      type_cast_1581_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1597_inst
    process(input_dim2x_x1_1517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_1517, tmp_var);
      type_cast_1597_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1634_inst
    process(inc_1631) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1631, tmp_var);
      type_cast_1634_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1660_inst
    process(inc72x_xinput_dim0x_x2_1650) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc72x_xinput_dim0x_x2_1650, tmp_var);
      type_cast_1660_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_1292_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1292_load_0_req_0;
      LOAD_padding_1292_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1292_load_0_req_1;
      LOAD_padding_1292_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1292_word_address_0;
      LOAD_padding_1292_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1364_load_0 ptr_deref_1263_load_0 ptr_deref_1251_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1364_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1263_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1251_load_0_req_0;
      ptr_deref_1364_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1263_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1251_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1364_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1263_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1251_load_0_req_1;
      ptr_deref_1364_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1263_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1251_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1364_word_address_0 & ptr_deref_1263_word_address_0 & ptr_deref_1251_word_address_0;
      ptr_deref_1364_data_0 <= data_out(95 downto 64);
      ptr_deref_1263_data_0 <= data_out(63 downto 32);
      ptr_deref_1251_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1306_load_0 ptr_deref_1273_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1306_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1273_load_0_req_0;
      ptr_deref_1306_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1273_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1306_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1273_load_0_req_1;
      ptr_deref_1306_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1273_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1306_word_address_0 & ptr_deref_1273_word_address_0;
      ptr_deref_1306_data_0 <= data_out(31 downto 16);
      ptr_deref_1273_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1322_load_0 ptr_deref_1289_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1322_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1289_load_0_req_0;
      ptr_deref_1322_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1289_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1322_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1289_load_0_req_1;
      ptr_deref_1322_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1289_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1322_word_address_0 & ptr_deref_1289_word_address_0;
      ptr_deref_1322_data_0 <= data_out(63 downto 32);
      ptr_deref_1289_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1334_load_0 ptr_deref_1346_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1334_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1346_load_0_req_0;
      ptr_deref_1334_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1346_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1334_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1346_load_0_req_1;
      ptr_deref_1334_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1346_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1334_word_address_0 & ptr_deref_1346_word_address_0;
      ptr_deref_1334_data_0 <= data_out(63 downto 32);
      ptr_deref_1346_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_1562_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1562_load_0_req_0;
      ptr_deref_1562_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1562_load_0_req_1;
      ptr_deref_1562_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1562_word_address_0;
      ptr_deref_1562_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_1592_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1592_store_0_req_0;
      ptr_deref_1592_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1592_store_0_req_1;
      ptr_deref_1592_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1592_word_address_0;
      data_in <= ptr_deref_1592_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1238_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_start_1238_inst_req_0;
      RPIPE_Block0_start_1238_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_start_1238_inst_req_1;
      RPIPE_Block0_start_1238_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1239 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1676_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1676_inst_req_0;
      WPIPE_Block0_done_1676_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1676_inst_req_1;
      WPIPE_Block0_done_1676_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1239;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4819_start: Boolean;
  signal convTransposeB_CP_4819_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_1686_inst_ack_1 : boolean;
  signal ptr_deref_1699_load_0_ack_1 : boolean;
  signal ptr_deref_1721_load_0_req_1 : boolean;
  signal ptr_deref_1721_load_0_ack_0 : boolean;
  signal RPIPE_Block1_start_1686_inst_req_1 : boolean;
  signal ptr_deref_1731_load_0_req_0 : boolean;
  signal ptr_deref_1731_load_0_ack_0 : boolean;
  signal RPIPE_Block1_start_1686_inst_req_0 : boolean;
  signal type_cast_1709_inst_req_0 : boolean;
  signal ptr_deref_1721_load_0_ack_1 : boolean;
  signal ptr_deref_1731_load_0_req_1 : boolean;
  signal type_cast_1735_inst_req_0 : boolean;
  signal type_cast_2132_inst_req_0 : boolean;
  signal type_cast_1735_inst_ack_0 : boolean;
  signal type_cast_2112_inst_ack_0 : boolean;
  signal type_cast_1709_inst_req_1 : boolean;
  signal ptr_deref_1699_load_0_ack_0 : boolean;
  signal RPIPE_Block1_start_1686_inst_ack_0 : boolean;
  signal type_cast_1709_inst_ack_0 : boolean;
  signal ptr_deref_1699_load_0_req_0 : boolean;
  signal ptr_deref_1699_load_0_req_1 : boolean;
  signal type_cast_1735_inst_req_1 : boolean;
  signal type_cast_1709_inst_ack_1 : boolean;
  signal type_cast_1735_inst_ack_1 : boolean;
  signal ptr_deref_1731_load_0_ack_1 : boolean;
  signal ptr_deref_1721_load_0_req_0 : boolean;
  signal type_cast_2132_inst_ack_0 : boolean;
  signal phi_stmt_1832_ack_0 : boolean;
  signal type_cast_2127_inst_req_0 : boolean;
  signal type_cast_2132_inst_req_1 : boolean;
  signal type_cast_2125_inst_ack_1 : boolean;
  signal type_cast_2132_inst_ack_1 : boolean;
  signal phi_stmt_2122_req_0 : boolean;
  signal type_cast_2125_inst_ack_0 : boolean;
  signal type_cast_1838_inst_req_1 : boolean;
  signal type_cast_2125_inst_req_1 : boolean;
  signal type_cast_2125_inst_req_0 : boolean;
  signal type_cast_2112_inst_req_1 : boolean;
  signal type_cast_2127_inst_ack_0 : boolean;
  signal type_cast_1957_inst_req_0 : boolean;
  signal type_cast_2112_inst_ack_1 : boolean;
  signal type_cast_1957_inst_ack_0 : boolean;
  signal ptr_deref_1747_load_0_req_0 : boolean;
  signal ptr_deref_1747_load_0_ack_0 : boolean;
  signal ptr_deref_1747_load_0_req_1 : boolean;
  signal ptr_deref_1747_load_0_ack_1 : boolean;
  signal if_stmt_2139_branch_ack_0 : boolean;
  signal LOAD_padding_1750_load_0_req_0 : boolean;
  signal LOAD_padding_1750_load_0_ack_0 : boolean;
  signal LOAD_padding_1750_load_0_req_1 : boolean;
  signal LOAD_padding_1750_load_0_ack_1 : boolean;
  signal type_cast_1754_inst_req_0 : boolean;
  signal type_cast_1754_inst_ack_0 : boolean;
  signal type_cast_1754_inst_req_1 : boolean;
  signal type_cast_1754_inst_ack_1 : boolean;
  signal ptr_deref_1764_load_0_req_0 : boolean;
  signal ptr_deref_1764_load_0_ack_0 : boolean;
  signal ptr_deref_1764_load_0_req_1 : boolean;
  signal ptr_deref_1764_load_0_ack_1 : boolean;
  signal type_cast_1768_inst_req_0 : boolean;
  signal type_cast_1768_inst_ack_0 : boolean;
  signal type_cast_1768_inst_req_1 : boolean;
  signal type_cast_1768_inst_ack_1 : boolean;
  signal ptr_deref_1780_load_0_req_0 : boolean;
  signal ptr_deref_1780_load_0_ack_0 : boolean;
  signal ptr_deref_1780_load_0_req_1 : boolean;
  signal ptr_deref_1780_load_0_ack_1 : boolean;
  signal ptr_deref_1792_load_0_req_0 : boolean;
  signal ptr_deref_1792_load_0_ack_0 : boolean;
  signal ptr_deref_1792_load_0_req_1 : boolean;
  signal ptr_deref_1792_load_0_ack_1 : boolean;
  signal ptr_deref_1804_load_0_req_0 : boolean;
  signal ptr_deref_1804_load_0_ack_0 : boolean;
  signal ptr_deref_1804_load_0_req_1 : boolean;
  signal ptr_deref_1804_load_0_ack_1 : boolean;
  signal type_cast_2112_inst_req_0 : boolean;
  signal phi_stmt_1826_ack_0 : boolean;
  signal phi_stmt_1826_req_0 : boolean;
  signal type_cast_1838_inst_ack_0 : boolean;
  signal if_stmt_2139_branch_ack_1 : boolean;
  signal ptr_deref_1816_load_0_req_0 : boolean;
  signal type_cast_1829_inst_ack_1 : boolean;
  signal ptr_deref_1816_load_0_ack_0 : boolean;
  signal type_cast_1838_inst_req_0 : boolean;
  signal ptr_deref_1816_load_0_req_1 : boolean;
  signal type_cast_1829_inst_req_1 : boolean;
  signal ptr_deref_1816_load_0_ack_1 : boolean;
  signal type_cast_1843_inst_req_0 : boolean;
  signal phi_stmt_1826_req_1 : boolean;
  signal type_cast_1843_inst_ack_0 : boolean;
  signal type_cast_1843_inst_req_1 : boolean;
  signal type_cast_1831_inst_ack_1 : boolean;
  signal type_cast_1843_inst_ack_1 : boolean;
  signal phi_stmt_2116_req_0 : boolean;
  signal type_cast_2119_inst_ack_1 : boolean;
  signal type_cast_1829_inst_ack_0 : boolean;
  signal type_cast_1848_inst_req_0 : boolean;
  signal type_cast_1831_inst_req_1 : boolean;
  signal type_cast_1848_inst_ack_0 : boolean;
  signal type_cast_1848_inst_req_1 : boolean;
  signal type_cast_1848_inst_ack_1 : boolean;
  signal type_cast_2119_inst_req_1 : boolean;
  signal phi_stmt_2122_ack_0 : boolean;
  signal type_cast_1829_inst_req_0 : boolean;
  signal phi_stmt_1954_ack_0 : boolean;
  signal type_cast_1970_inst_req_0 : boolean;
  signal type_cast_1970_inst_ack_0 : boolean;
  signal type_cast_1970_inst_req_1 : boolean;
  signal type_cast_1831_inst_ack_0 : boolean;
  signal type_cast_1970_inst_ack_1 : boolean;
  signal phi_stmt_2116_ack_0 : boolean;
  signal type_cast_2119_inst_ack_0 : boolean;
  signal phi_stmt_2116_req_1 : boolean;
  signal type_cast_2000_inst_req_0 : boolean;
  signal type_cast_1831_inst_req_0 : boolean;
  signal type_cast_2000_inst_ack_0 : boolean;
  signal type_cast_2121_inst_ack_1 : boolean;
  signal type_cast_2000_inst_req_1 : boolean;
  signal type_cast_2000_inst_ack_1 : boolean;
  signal type_cast_2119_inst_req_0 : boolean;
  signal phi_stmt_1954_req_1 : boolean;
  signal type_cast_2121_inst_req_1 : boolean;
  signal if_stmt_2091_branch_ack_0 : boolean;
  signal phi_stmt_2122_req_1 : boolean;
  signal array_obj_ref_2006_index_offset_req_0 : boolean;
  signal array_obj_ref_2006_index_offset_ack_0 : boolean;
  signal array_obj_ref_2006_index_offset_req_1 : boolean;
  signal array_obj_ref_2006_index_offset_ack_1 : boolean;
  signal type_cast_2127_inst_ack_1 : boolean;
  signal type_cast_2127_inst_req_1 : boolean;
  signal addr_of_2007_final_reg_req_0 : boolean;
  signal addr_of_2007_final_reg_ack_0 : boolean;
  signal addr_of_2007_final_reg_req_1 : boolean;
  signal addr_of_2007_final_reg_ack_1 : boolean;
  signal phi_stmt_1954_req_0 : boolean;
  signal phi_stmt_1832_req_0 : boolean;
  signal if_stmt_2139_branch_req_0 : boolean;
  signal ptr_deref_2011_load_0_req_0 : boolean;
  signal ptr_deref_2011_load_0_ack_0 : boolean;
  signal ptr_deref_2011_load_0_req_1 : boolean;
  signal ptr_deref_2011_load_0_ack_1 : boolean;
  signal type_cast_2121_inst_ack_0 : boolean;
  signal type_cast_1957_inst_ack_1 : boolean;
  signal WPIPE_Block1_done_2147_inst_ack_1 : boolean;
  signal type_cast_2121_inst_req_0 : boolean;
  signal type_cast_2031_inst_req_0 : boolean;
  signal phi_stmt_1832_req_1 : boolean;
  signal type_cast_2031_inst_ack_0 : boolean;
  signal if_stmt_2091_branch_ack_1 : boolean;
  signal type_cast_2031_inst_req_1 : boolean;
  signal type_cast_1838_inst_ack_1 : boolean;
  signal type_cast_2031_inst_ack_1 : boolean;
  signal type_cast_1957_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2147_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2147_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2147_inst_req_0 : boolean;
  signal array_obj_ref_2037_index_offset_req_0 : boolean;
  signal array_obj_ref_2037_index_offset_ack_0 : boolean;
  signal array_obj_ref_2037_index_offset_req_1 : boolean;
  signal array_obj_ref_2037_index_offset_ack_1 : boolean;
  signal addr_of_2038_final_reg_req_0 : boolean;
  signal addr_of_2038_final_reg_ack_0 : boolean;
  signal addr_of_2038_final_reg_req_1 : boolean;
  signal addr_of_2038_final_reg_ack_1 : boolean;
  signal ptr_deref_2041_store_0_req_0 : boolean;
  signal ptr_deref_2041_store_0_ack_0 : boolean;
  signal ptr_deref_2041_store_0_req_1 : boolean;
  signal ptr_deref_2041_store_0_ack_1 : boolean;
  signal type_cast_2047_inst_req_0 : boolean;
  signal type_cast_2047_inst_ack_0 : boolean;
  signal type_cast_2047_inst_req_1 : boolean;
  signal type_cast_2047_inst_ack_1 : boolean;
  signal if_stmt_2060_branch_req_0 : boolean;
  signal if_stmt_2060_branch_ack_1 : boolean;
  signal if_stmt_2060_branch_ack_0 : boolean;
  signal type_cast_2084_inst_req_0 : boolean;
  signal type_cast_2084_inst_ack_0 : boolean;
  signal type_cast_2084_inst_req_1 : boolean;
  signal type_cast_2084_inst_ack_1 : boolean;
  signal if_stmt_2091_branch_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4819_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4819_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4819_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4819_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4819: Block -- control-path 
    signal convTransposeB_CP_4819_elements: BooleanArray(112 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4819_elements(0) <= convTransposeB_CP_4819_start;
    convTransposeB_CP_4819_symbol <= convTransposeB_CP_4819_elements(72);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1684/assign_stmt_1687/RPIPE_Block1_start_1686_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1684/assign_stmt_1687/RPIPE_Block1_start_1686_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1684/$entry
      -- CP-element group 0: 	 branch_block_stmt_1684/branch_block_stmt_1684__entry__
      -- CP-element group 0: 	 branch_block_stmt_1684/assign_stmt_1687__entry__
      -- CP-element group 0: 	 branch_block_stmt_1684/assign_stmt_1687/$entry
      -- CP-element group 0: 	 branch_block_stmt_1684/assign_stmt_1687/RPIPE_Block1_start_1686_sample_start_
      -- 
    rr_4877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(0), ack => RPIPE_Block1_start_1686_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1684/assign_stmt_1687/RPIPE_Block1_start_1686_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1684/assign_stmt_1687/RPIPE_Block1_start_1686_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1684/assign_stmt_1687/RPIPE_Block1_start_1686_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1684/assign_stmt_1687/RPIPE_Block1_start_1686_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1684/assign_stmt_1687/RPIPE_Block1_start_1686_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1684/assign_stmt_1687/RPIPE_Block1_start_1686_update_start_
      -- 
    ra_4878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1686_inst_ack_0, ack => convTransposeB_CP_4819_elements(1)); -- 
    cr_4882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(1), ack => RPIPE_Block1_start_1686_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	12 
    -- CP-element group 2:  members (265) 
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1687/RPIPE_Block1_start_1686_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1687/RPIPE_Block1_start_1686_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1709_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1709_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1735_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1735_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1709_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1735_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1687__exit__
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823__entry__
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1687/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1687/RPIPE_Block1_start_1686_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1754_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1754_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1754_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1768_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1768_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1768_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Update/word_access_complete/word_0/cr
      -- 
    ca_4883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1686_inst_ack_1, ack => convTransposeB_CP_4819_elements(2)); -- 
    cr_4994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1721_load_0_req_1); -- 
    rr_5033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1731_load_0_req_0); -- 
    cr_5044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1731_load_0_req_1); -- 
    cr_4949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => type_cast_1709_inst_req_1); -- 
    rr_4919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1699_load_0_req_0); -- 
    cr_4930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1699_load_0_req_1); -- 
    cr_5063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => type_cast_1735_inst_req_1); -- 
    rr_4983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1721_load_0_req_0); -- 
    rr_5097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1747_load_0_req_0); -- 
    cr_5108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1747_load_0_req_1); -- 
    rr_5130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => LOAD_padding_1750_load_0_req_0); -- 
    cr_5141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => LOAD_padding_1750_load_0_req_1); -- 
    cr_5160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => type_cast_1754_inst_req_1); -- 
    rr_5194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1764_load_0_req_0); -- 
    cr_5205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1764_load_0_req_1); -- 
    cr_5224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => type_cast_1768_inst_req_1); -- 
    rr_5258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1780_load_0_req_0); -- 
    cr_5269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1780_load_0_req_1); -- 
    rr_5308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1792_load_0_req_0); -- 
    cr_5319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1792_load_0_req_1); -- 
    rr_5358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1804_load_0_req_0); -- 
    cr_5369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1804_load_0_req_1); -- 
    rr_5408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1816_load_0_req_0); -- 
    cr_5419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(2), ack => ptr_deref_1816_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Sample/$exit
      -- 
    ra_4920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1699_load_0_ack_0, ack => convTransposeB_CP_4819_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Update/ptr_deref_1699_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1709_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Update/ptr_deref_1699_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Update/ptr_deref_1699_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1709_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1699_Update/ptr_deref_1699_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1709_Sample/$entry
      -- 
    ca_4931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1699_load_0_ack_1, ack => convTransposeB_CP_4819_elements(4)); -- 
    rr_4944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(4), ack => type_cast_1709_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1709_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1709_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1709_Sample/ra
      -- 
    ra_4945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1709_inst_ack_0, ack => convTransposeB_CP_4819_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	31 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1709_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1709_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1709_Update/ca
      -- 
    ca_4950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1709_inst_ack_1, ack => convTransposeB_CP_4819_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Sample/word_access_start/word_0/$exit
      -- 
    ra_4984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1721_load_0_ack_0, ack => convTransposeB_CP_4819_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	31 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Update/ptr_deref_1721_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Update/ptr_deref_1721_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Update/ptr_deref_1721_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Update/ptr_deref_1721_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1721_Update/word_access_complete/word_0/$exit
      -- 
    ca_4995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1721_load_0_ack_1, ack => convTransposeB_CP_4819_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Sample/word_access_start/word_0/ra
      -- CP-element group 9: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_sample_completed_
      -- 
    ra_5034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1731_load_0_ack_0, ack => convTransposeB_CP_4819_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (12) 
      -- CP-element group 10: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1735_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Update/ptr_deref_1731_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Update/ptr_deref_1731_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Update/ptr_deref_1731_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1735_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1735_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Update/ptr_deref_1731_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1731_Update/word_access_complete/word_0/$exit
      -- 
    ca_5045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1731_load_0_ack_1, ack => convTransposeB_CP_4819_elements(10)); -- 
    rr_5058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(10), ack => type_cast_1735_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1735_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1735_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1735_Sample/ra
      -- 
    ra_5059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1735_inst_ack_0, ack => convTransposeB_CP_4819_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	31 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1735_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1735_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1735_Update/ca
      -- 
    ca_5064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1735_inst_ack_1, ack => convTransposeB_CP_4819_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Sample/word_access_start/word_0/ra
      -- 
    ra_5098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1747_load_0_ack_0, ack => convTransposeB_CP_4819_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	31 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Update/ptr_deref_1747_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Update/ptr_deref_1747_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Update/ptr_deref_1747_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1747_Update/ptr_deref_1747_Merge/merge_ack
      -- 
    ca_5109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1747_load_0_ack_1, ack => convTransposeB_CP_4819_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Sample/word_access_start/word_0/ra
      -- 
    ra_5131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1750_load_0_ack_0, ack => convTransposeB_CP_4819_elements(15)); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (12) 
      -- CP-element group 16: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Update/LOAD_padding_1750_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Update/LOAD_padding_1750_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Update/LOAD_padding_1750_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/LOAD_padding_1750_Update/LOAD_padding_1750_Merge/merge_ack
      -- CP-element group 16: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1754_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1754_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1754_Sample/rr
      -- 
    ca_5142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1750_load_0_ack_1, ack => convTransposeB_CP_4819_elements(16)); -- 
    rr_5155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(16), ack => type_cast_1754_inst_req_0); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1754_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1754_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1754_Sample/ra
      -- 
    ra_5156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1754_inst_ack_0, ack => convTransposeB_CP_4819_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	31 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1754_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1754_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1754_Update/ca
      -- 
    ca_5161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1754_inst_ack_1, ack => convTransposeB_CP_4819_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Sample/word_access_start/word_0/ra
      -- 
    ra_5195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1764_load_0_ack_0, ack => convTransposeB_CP_4819_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (12) 
      -- CP-element group 20: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Update/ptr_deref_1764_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Update/ptr_deref_1764_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Update/ptr_deref_1764_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1764_Update/ptr_deref_1764_Merge/merge_ack
      -- CP-element group 20: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1768_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1768_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1768_Sample/rr
      -- 
    ca_5206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1764_load_0_ack_1, ack => convTransposeB_CP_4819_elements(20)); -- 
    rr_5219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(20), ack => type_cast_1768_inst_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1768_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1768_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1768_Sample/ra
      -- 
    ra_5220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1768_inst_ack_0, ack => convTransposeB_CP_4819_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	31 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1768_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1768_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/type_cast_1768_Update/ca
      -- 
    ca_5225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1768_inst_ack_1, ack => convTransposeB_CP_4819_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Sample/word_access_start/word_0/ra
      -- 
    ra_5259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1780_load_0_ack_0, ack => convTransposeB_CP_4819_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	31 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Update/ptr_deref_1780_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Update/ptr_deref_1780_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Update/ptr_deref_1780_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1780_Update/ptr_deref_1780_Merge/merge_ack
      -- 
    ca_5270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1780_load_0_ack_1, ack => convTransposeB_CP_4819_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Sample/word_access_start/word_0/ra
      -- 
    ra_5309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1792_load_0_ack_0, ack => convTransposeB_CP_4819_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Update/ptr_deref_1792_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Update/ptr_deref_1792_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Update/ptr_deref_1792_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1792_Update/ptr_deref_1792_Merge/merge_ack
      -- 
    ca_5320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1792_load_0_ack_1, ack => convTransposeB_CP_4819_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Sample/word_access_start/word_0/ra
      -- 
    ra_5359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1804_load_0_ack_0, ack => convTransposeB_CP_4819_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Update/ptr_deref_1804_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Update/ptr_deref_1804_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Update/ptr_deref_1804_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1804_Update/ptr_deref_1804_Merge/merge_ack
      -- 
    ca_5370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1804_load_0_ack_1, ack => convTransposeB_CP_4819_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Sample/word_access_start/word_0/ra
      -- 
    ra_5409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1816_load_0_ack_0, ack => convTransposeB_CP_4819_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Update/ptr_deref_1816_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Update/ptr_deref_1816_Merge/$exit
      -- CP-element group 30: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Update/ptr_deref_1816_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/ptr_deref_1816_Update/ptr_deref_1816_Merge/merge_ack
      -- 
    ca_5420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1816_load_0_ack_1, ack => convTransposeB_CP_4819_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	22 
    -- CP-element group 31: 	24 
    -- CP-element group 31: 	14 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	18 
    -- CP-element group 31: 	6 
    -- CP-element group 31: 	8 
    -- CP-element group 31: 	12 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	73 
    -- CP-element group 31: 	74 
    -- CP-element group 31: 	75 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823/$exit
      -- CP-element group 31: 	 branch_block_stmt_1684/assign_stmt_1696_to_assign_stmt_1823__exit__
      -- CP-element group 31: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1829/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1829/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1829/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1829/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1829/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1829/$entry
      -- CP-element group 31: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/$entry
      -- CP-element group 31: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/$entry
      -- CP-element group 31: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- 
    cr_5867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(31), ack => type_cast_1829_inst_req_1); -- 
    rr_5862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(31), ack => type_cast_1829_inst_req_0); -- 
    convTransposeB_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(22) & convTransposeB_CP_4819_elements(24) & convTransposeB_CP_4819_elements(14) & convTransposeB_CP_4819_elements(26) & convTransposeB_CP_4819_elements(28) & convTransposeB_CP_4819_elements(30) & convTransposeB_CP_4819_elements(18) & convTransposeB_CP_4819_elements(6) & convTransposeB_CP_4819_elements(8) & convTransposeB_CP_4819_elements(12);
      gj_convTransposeB_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	88 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1843_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1843_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1843_Sample/ra
      -- 
    ra_5437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1843_inst_ack_0, ack => convTransposeB_CP_4819_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	88 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1843_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1843_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1843_Update/ca
      -- 
    ca_5442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1843_inst_ack_1, ack => convTransposeB_CP_4819_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	88 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1848_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1848_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1848_Sample/ra
      -- 
    ra_5451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1848_inst_ack_0, ack => convTransposeB_CP_4819_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	88 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1848_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1848_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1848_Update/ca
      -- 
    ca_5456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1848_inst_ack_1, ack => convTransposeB_CP_4819_elements(35)); -- 
    -- CP-element group 36:  join  transition  place  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	33 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	92 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951__exit__
      -- CP-element group 36: 	 branch_block_stmt_1684/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 36: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/$exit
      -- CP-element group 36: 	 branch_block_stmt_1684/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/$entry
      -- CP-element group 36: 	 branch_block_stmt_1684/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1954/$entry
      -- CP-element group 36: 	 branch_block_stmt_1684/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- 
    convTransposeB_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(33) & convTransposeB_CP_4819_elements(35);
      gj_convTransposeB_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	94 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_1970_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_1970_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_1970_Sample/ra
      -- 
    ra_5468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1970_inst_ack_0, ack => convTransposeB_CP_4819_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	94 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	47 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_1970_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_1970_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_1970_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2000_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2000_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2000_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2031_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2031_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2031_Sample/rr
      -- 
    ca_5473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1970_inst_ack_1, ack => convTransposeB_CP_4819_elements(38)); -- 
    rr_5591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(38), ack => type_cast_2031_inst_req_0); -- 
    rr_5481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(38), ack => type_cast_2000_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2000_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2000_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2000_Sample/ra
      -- 
    ra_5482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2000_inst_ack_0, ack => convTransposeB_CP_4819_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	94 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (16) 
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2000_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2000_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2000_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_index_resized_1
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_index_scaled_1
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_index_computed_1
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_index_resize_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_index_resize_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_index_resize_1/index_resize_req
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_index_resize_1/index_resize_ack
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_index_scale_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_index_scale_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_index_scale_1/scale_rename_req
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_index_scale_1/scale_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_final_index_sum_regn_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_final_index_sum_regn_Sample/req
      -- 
    ca_5487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2000_inst_ack_1, ack => convTransposeB_CP_4819_elements(40)); -- 
    req_5512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(40), ack => array_obj_ref_2006_index_offset_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_final_index_sum_regn_sample_complete
      -- CP-element group 41: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_final_index_sum_regn_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_final_index_sum_regn_Sample/ack
      -- 
    ack_5513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2006_index_offset_ack_0, ack => convTransposeB_CP_4819_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	94 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (11) 
      -- CP-element group 42: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2007_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_offset_calculated
      -- CP-element group 42: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_final_index_sum_regn_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_final_index_sum_regn_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2007_request/$entry
      -- CP-element group 42: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2007_request/req
      -- 
    ack_5518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2006_index_offset_ack_1, ack => convTransposeB_CP_4819_elements(42)); -- 
    req_5527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(42), ack => addr_of_2007_final_reg_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2007_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2007_request/$exit
      -- CP-element group 43: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2007_request/ack
      -- 
    ack_5528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2007_final_reg_ack_0, ack => convTransposeB_CP_4819_elements(43)); -- 
    -- CP-element group 44:  join  fork  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	94 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (24) 
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2007_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2007_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2007_complete/ack
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_base_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_word_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_base_address_resized
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_base_addr_resize/$entry
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_base_addr_resize/$exit
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_base_addr_resize/base_resize_req
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_base_addr_resize/base_resize_ack
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_word_addrgen/$entry
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_word_addrgen/$exit
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_word_addrgen/root_register_req
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_word_addrgen/root_register_ack
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Sample/word_access_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Sample/word_access_start/word_0/rr
      -- 
    ack_5533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2007_final_reg_ack_1, ack => convTransposeB_CP_4819_elements(44)); -- 
    rr_5566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(44), ack => ptr_deref_2011_load_0_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Sample/word_access_start/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Sample/word_access_start/word_0/ra
      -- 
    ra_5567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_load_0_ack_0, ack => convTransposeB_CP_4819_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	94 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	53 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Update/word_access_complete/word_0/ca
      -- CP-element group 46: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Update/ptr_deref_2011_Merge/$entry
      -- CP-element group 46: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Update/ptr_deref_2011_Merge/$exit
      -- CP-element group 46: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Update/ptr_deref_2011_Merge/merge_req
      -- CP-element group 46: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Update/ptr_deref_2011_Merge/merge_ack
      -- 
    ca_5578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_load_0_ack_1, ack => convTransposeB_CP_4819_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	38 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2031_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2031_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2031_Sample/ra
      -- 
    ra_5592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2031_inst_ack_0, ack => convTransposeB_CP_4819_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	94 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (16) 
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2031_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2031_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2031_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_index_resized_1
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_index_scaled_1
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_index_computed_1
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_index_resize_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_index_resize_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_index_resize_1/index_resize_req
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_index_resize_1/index_resize_ack
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_index_scale_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_index_scale_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_index_scale_1/scale_rename_req
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_index_scale_1/scale_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_final_index_sum_regn_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_final_index_sum_regn_Sample/req
      -- 
    ca_5597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2031_inst_ack_1, ack => convTransposeB_CP_4819_elements(48)); -- 
    req_5622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(48), ack => array_obj_ref_2037_index_offset_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_final_index_sum_regn_sample_complete
      -- CP-element group 49: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_final_index_sum_regn_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_final_index_sum_regn_Sample/ack
      -- 
    ack_5623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2037_index_offset_ack_0, ack => convTransposeB_CP_4819_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	94 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (11) 
      -- CP-element group 50: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2038_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_offset_calculated
      -- CP-element group 50: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_final_index_sum_regn_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_final_index_sum_regn_Update/ack
      -- CP-element group 50: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2038_request/$entry
      -- CP-element group 50: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2038_request/req
      -- 
    ack_5628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2037_index_offset_ack_1, ack => convTransposeB_CP_4819_elements(50)); -- 
    req_5637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(50), ack => addr_of_2038_final_reg_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2038_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2038_request/$exit
      -- CP-element group 51: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2038_request/ack
      -- 
    ack_5638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2038_final_reg_ack_0, ack => convTransposeB_CP_4819_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	94 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (19) 
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2038_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2038_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2038_complete/ack
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_word_addrgen/root_register_ack
      -- 
    ack_5643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2038_final_reg_ack_1, ack => convTransposeB_CP_4819_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	46 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Sample/ptr_deref_2041_Split/$entry
      -- CP-element group 53: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Sample/ptr_deref_2041_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Sample/ptr_deref_2041_Split/split_req
      -- CP-element group 53: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Sample/ptr_deref_2041_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Sample/word_access_start/word_0/rr
      -- 
    rr_5681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(53), ack => ptr_deref_2041_store_0_req_0); -- 
    convTransposeB_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(46) & convTransposeB_CP_4819_elements(52);
      gj_convTransposeB_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Sample/word_access_start/word_0/ra
      -- 
    ra_5682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2041_store_0_ack_0, ack => convTransposeB_CP_4819_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	94 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Update/word_access_complete/word_0/ca
      -- 
    ca_5693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2041_store_0_ack_1, ack => convTransposeB_CP_4819_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	94 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2047_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2047_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2047_Sample/ra
      -- 
    ra_5702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2047_inst_ack_0, ack => convTransposeB_CP_4819_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	94 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2047_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2047_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2047_Update/ca
      -- 
    ca_5707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2047_inst_ack_1, ack => convTransposeB_CP_4819_elements(57)); -- 
    -- CP-element group 58:  branch  join  transition  place  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	49 
    -- CP-element group 58: 	55 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (10) 
      -- CP-element group 58: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059__exit__
      -- CP-element group 58: 	 branch_block_stmt_1684/if_stmt_2060__entry__
      -- CP-element group 58: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/$exit
      -- CP-element group 58: 	 branch_block_stmt_1684/if_stmt_2060_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1684/if_stmt_2060_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_1684/if_stmt_2060_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_1684/if_stmt_2060_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_1684/R_cmp_2061_place
      -- CP-element group 58: 	 branch_block_stmt_1684/if_stmt_2060_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1684/if_stmt_2060_else_link/$entry
      -- 
    branch_req_5715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(58), ack => if_stmt_2060_branch_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(41) & convTransposeB_CP_4819_elements(49) & convTransposeB_CP_4819_elements(55) & convTransposeB_CP_4819_elements(57);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	89 
    -- CP-element group 59: 	90 
    -- CP-element group 59:  members (24) 
      -- CP-element group 59: 	 branch_block_stmt_1684/merge_stmt_2066_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/$entry
      -- CP-element group 59: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/$entry
      -- CP-element group 59: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1684/merge_stmt_2066__exit__
      -- CP-element group 59: 	 branch_block_stmt_1684/assign_stmt_2072__entry__
      -- CP-element group 59: 	 branch_block_stmt_1684/assign_stmt_2072__exit__
      -- CP-element group 59: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody
      -- CP-element group 59: 	 branch_block_stmt_1684/merge_stmt_2066_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_1684/merge_stmt_2066_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1684/merge_stmt_2066_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1684/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_1684/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Update/cr
      -- CP-element group 59: 	 branch_block_stmt_1684/if_stmt_2060_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1684/if_stmt_2060_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1684/whilex_xbody_ifx_xthen
      -- CP-element group 59: 	 branch_block_stmt_1684/assign_stmt_2072/$entry
      -- CP-element group 59: 	 branch_block_stmt_1684/assign_stmt_2072/$exit
      -- 
    if_choice_transition_5720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2060_branch_ack_1, ack => convTransposeB_CP_4819_elements(59)); -- 
    rr_5943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(59), ack => type_cast_1957_inst_req_0); -- 
    cr_5948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(59), ack => type_cast_1957_inst_req_1); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (18) 
      -- CP-element group 60: 	 branch_block_stmt_1684/merge_stmt_2074_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_1684/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_1684/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_1684/merge_stmt_2074_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_1684/merge_stmt_2074_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_1684/merge_stmt_2074_PhiAck/dummy
      -- CP-element group 60: 	 branch_block_stmt_1684/merge_stmt_2074__exit__
      -- CP-element group 60: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090__entry__
      -- CP-element group 60: 	 branch_block_stmt_1684/if_stmt_2060_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_1684/if_stmt_2060_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_1684/whilex_xbody_ifx_xelse
      -- CP-element group 60: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/$entry
      -- CP-element group 60: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/type_cast_2084_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/type_cast_2084_update_start_
      -- CP-element group 60: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/type_cast_2084_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/type_cast_2084_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/type_cast_2084_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/type_cast_2084_Update/cr
      -- 
    else_choice_transition_5724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2060_branch_ack_0, ack => convTransposeB_CP_4819_elements(60)); -- 
    rr_5740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(60), ack => type_cast_2084_inst_req_0); -- 
    cr_5745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(60), ack => type_cast_2084_inst_req_1); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/type_cast_2084_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/type_cast_2084_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/type_cast_2084_Sample/ra
      -- 
    ra_5741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2084_inst_ack_0, ack => convTransposeB_CP_4819_elements(61)); -- 
    -- CP-element group 62:  branch  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (13) 
      -- CP-element group 62: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090__exit__
      -- CP-element group 62: 	 branch_block_stmt_1684/if_stmt_2091__entry__
      -- CP-element group 62: 	 branch_block_stmt_1684/if_stmt_2091_else_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_1684/if_stmt_2091_if_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/$exit
      -- CP-element group 62: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/type_cast_2084_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/type_cast_2084_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1684/assign_stmt_2080_to_assign_stmt_2090/type_cast_2084_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1684/if_stmt_2091_dead_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_1684/if_stmt_2091_eval_test/$entry
      -- CP-element group 62: 	 branch_block_stmt_1684/if_stmt_2091_eval_test/$exit
      -- CP-element group 62: 	 branch_block_stmt_1684/if_stmt_2091_eval_test/branch_req
      -- CP-element group 62: 	 branch_block_stmt_1684/R_cmp77_2092_place
      -- 
    ca_5746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2084_inst_ack_1, ack => convTransposeB_CP_4819_elements(62)); -- 
    branch_req_5754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(62), ack => if_stmt_2091_branch_req_0); -- 
    -- CP-element group 63:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (18) 
      -- CP-element group 63: 	 branch_block_stmt_1684/merge_stmt_2097_PhiReqMerge
      -- CP-element group 63: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/type_cast_2112_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_1684/ifx_xelse_ifx_xthen79_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_1684/ifx_xelse_ifx_xthen79_PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_1684/merge_stmt_2097_PhiAck/$entry
      -- CP-element group 63: 	 branch_block_stmt_1684/merge_stmt_2097_PhiAck/$exit
      -- CP-element group 63: 	 branch_block_stmt_1684/merge_stmt_2097_PhiAck/dummy
      -- CP-element group 63: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/type_cast_2112_Update/cr
      -- CP-element group 63: 	 branch_block_stmt_1684/merge_stmt_2097__exit__
      -- CP-element group 63: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113__entry__
      -- CP-element group 63: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/type_cast_2112_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/type_cast_2112_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1684/ifx_xelse_ifx_xthen79
      -- CP-element group 63: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/$entry
      -- CP-element group 63: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/type_cast_2112_update_start_
      -- CP-element group 63: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/type_cast_2112_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1684/if_stmt_2091_if_link/if_choice_transition
      -- CP-element group 63: 	 branch_block_stmt_1684/if_stmt_2091_if_link/$exit
      -- 
    if_choice_transition_5759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2091_branch_ack_1, ack => convTransposeB_CP_4819_elements(63)); -- 
    cr_5781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(63), ack => type_cast_2112_inst_req_1); -- 
    rr_5776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(63), ack => type_cast_2112_inst_req_0); -- 
    -- CP-element group 64:  fork  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	95 
    -- CP-element group 64: 	96 
    -- CP-element group 64: 	98 
    -- CP-element group 64: 	99 
    -- CP-element group 64:  members (20) 
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2127/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2121/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2127/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2121/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2127/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2121/$entry
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2127/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2127/$entry
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/$entry
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2121/SplitProtocol/Update/cr
      -- CP-element group 64: 	 branch_block_stmt_1684/if_stmt_2091_else_link/else_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2127/SplitProtocol/Update/cr
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2121/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1684/if_stmt_2091_else_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/$entry
      -- CP-element group 64: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2121/SplitProtocol/Sample/rr
      -- 
    else_choice_transition_5763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2091_branch_ack_0, ack => convTransposeB_CP_4819_elements(64)); -- 
    rr_6040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(64), ack => type_cast_2127_inst_req_0); -- 
    cr_6022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(64), ack => type_cast_2121_inst_req_1); -- 
    cr_6045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(64), ack => type_cast_2127_inst_req_1); -- 
    rr_6017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(64), ack => type_cast_2121_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/type_cast_2112_Sample/ra
      -- CP-element group 65: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/type_cast_2112_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/type_cast_2112_sample_completed_
      -- 
    ra_5777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2112_inst_ack_0, ack => convTransposeB_CP_4819_elements(65)); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	102 
    -- CP-element group 66: 	103 
    -- CP-element group 66: 	105 
    -- CP-element group 66: 	106 
    -- CP-element group 66:  members (23) 
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/type_cast_2112_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2119/$entry
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2125/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2125/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2125/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2119/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2125/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2125/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/type_cast_2112_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2125/$entry
      -- CP-element group 66: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113__exit__
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend
      -- CP-element group 66: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/type_cast_2112_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/$entry
      -- CP-element group 66: 	 branch_block_stmt_1684/assign_stmt_2103_to_assign_stmt_2113/$exit
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/$entry
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2119/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2119/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2119/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2119/SplitProtocol/Sample/$entry
      -- 
    ca_5782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2112_inst_ack_1, ack => convTransposeB_CP_4819_elements(66)); -- 
    cr_6094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(66), ack => type_cast_2125_inst_req_1); -- 
    rr_6089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(66), ack => type_cast_2125_inst_req_0); -- 
    cr_6071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(66), ack => type_cast_2119_inst_req_1); -- 
    rr_6066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(66), ack => type_cast_2119_inst_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	112 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/type_cast_2132_Sample/ra
      -- CP-element group 67: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/type_cast_2132_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/type_cast_2132_sample_completed_
      -- 
    ra_5794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2132_inst_ack_0, ack => convTransposeB_CP_4819_elements(67)); -- 
    -- CP-element group 68:  branch  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	112 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (13) 
      -- CP-element group 68: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/type_cast_2132_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/type_cast_2132_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_1684/if_stmt_2139_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138__exit__
      -- CP-element group 68: 	 branch_block_stmt_1684/if_stmt_2139__entry__
      -- CP-element group 68: 	 branch_block_stmt_1684/if_stmt_2139_else_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1684/R_cmp89_2140_place
      -- CP-element group 68: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/type_cast_2132_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_1684/if_stmt_2139_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1684/if_stmt_2139_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1684/if_stmt_2139_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1684/if_stmt_2139_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/$exit
      -- 
    ca_5799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2132_inst_ack_1, ack => convTransposeB_CP_4819_elements(68)); -- 
    branch_req_5807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(68), ack => if_stmt_2139_branch_req_0); -- 
    -- CP-element group 69:  merge  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (15) 
      -- CP-element group 69: 	 branch_block_stmt_1684/merge_stmt_2145_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1684/assign_stmt_2149/$entry
      -- CP-element group 69: 	 branch_block_stmt_1684/ifx_xend_whilex_xend
      -- CP-element group 69: 	 branch_block_stmt_1684/assign_stmt_2149/WPIPE_Block1_done_2147_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_1684/merge_stmt_2145_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1684/merge_stmt_2145_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1684/ifx_xend_whilex_xend_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1684/merge_stmt_2145_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1684/merge_stmt_2145__exit__
      -- CP-element group 69: 	 branch_block_stmt_1684/assign_stmt_2149__entry__
      -- CP-element group 69: 	 branch_block_stmt_1684/if_stmt_2139_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1684/if_stmt_2139_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1684/ifx_xend_whilex_xend_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1684/assign_stmt_2149/WPIPE_Block1_done_2147_Sample/req
      -- CP-element group 69: 	 branch_block_stmt_1684/assign_stmt_2149/WPIPE_Block1_done_2147_Sample/$entry
      -- 
    if_choice_transition_5812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2139_branch_ack_1, ack => convTransposeB_CP_4819_elements(69)); -- 
    req_5829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(69), ack => WPIPE_Block1_done_2147_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	78 
    -- CP-element group 70: 	79 
    -- CP-element group 70: 	81 
    -- CP-element group 70: 	82 
    -- CP-element group 70:  members (20) 
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/type_cast_1838/SplitProtocol/Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/$entry
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/$entry
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/type_cast_1838/SplitProtocol/Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/type_cast_1838/$entry
      -- CP-element group 70: 	 branch_block_stmt_1684/if_stmt_2139_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1684/if_stmt_2139_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/type_cast_1838/SplitProtocol/Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1831/SplitProtocol/Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1831/SplitProtocol/Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1831/SplitProtocol/Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/type_cast_1838/SplitProtocol/Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1831/SplitProtocol/Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1831/SplitProtocol/$entry
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1831/$entry
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/type_cast_1838/SplitProtocol/$entry
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/$entry
      -- CP-element group 70: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/$entry
      -- 
    else_choice_transition_5816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2139_branch_ack_0, ack => convTransposeB_CP_4819_elements(70)); -- 
    cr_5893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(70), ack => type_cast_1838_inst_req_1); -- 
    rr_5888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(70), ack => type_cast_1838_inst_req_0); -- 
    cr_5916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(70), ack => type_cast_1831_inst_req_1); -- 
    rr_5911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(70), ack => type_cast_1831_inst_req_0); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_1684/assign_stmt_2149/WPIPE_Block1_done_2147_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1684/assign_stmt_2149/WPIPE_Block1_done_2147_Update/req
      -- CP-element group 71: 	 branch_block_stmt_1684/assign_stmt_2149/WPIPE_Block1_done_2147_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1684/assign_stmt_2149/WPIPE_Block1_done_2147_Sample/ack
      -- CP-element group 71: 	 branch_block_stmt_1684/assign_stmt_2149/WPIPE_Block1_done_2147_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1684/assign_stmt_2149/WPIPE_Block1_done_2147_update_start_
      -- 
    ack_5830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2147_inst_ack_0, ack => convTransposeB_CP_4819_elements(71)); -- 
    req_5834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(71), ack => WPIPE_Block1_done_2147_inst_req_1); -- 
    -- CP-element group 72:  transition  place  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (16) 
      -- CP-element group 72: 	 branch_block_stmt_1684/merge_stmt_2151_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_1684/assign_stmt_2149/$exit
      -- CP-element group 72: 	 branch_block_stmt_1684/return___PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_1684/return___PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_1684/merge_stmt_2151_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_1684/merge_stmt_2151_PhiAck/$exit
      -- CP-element group 72: 	 branch_block_stmt_1684/merge_stmt_2151_PhiAck/dummy
      -- CP-element group 72: 	 $exit
      -- CP-element group 72: 	 branch_block_stmt_1684/$exit
      -- CP-element group 72: 	 branch_block_stmt_1684/branch_block_stmt_1684__exit__
      -- CP-element group 72: 	 branch_block_stmt_1684/assign_stmt_2149__exit__
      -- CP-element group 72: 	 branch_block_stmt_1684/return__
      -- CP-element group 72: 	 branch_block_stmt_1684/merge_stmt_2151__exit__
      -- CP-element group 72: 	 branch_block_stmt_1684/assign_stmt_2149/WPIPE_Block1_done_2147_Update/ack
      -- CP-element group 72: 	 branch_block_stmt_1684/assign_stmt_2149/WPIPE_Block1_done_2147_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1684/assign_stmt_2149/WPIPE_Block1_done_2147_update_completed_
      -- 
    ack_5835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2147_inst_ack_1, ack => convTransposeB_CP_4819_elements(72)); -- 
    -- CP-element group 73:  transition  output  delay-element  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	31 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	77 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_req
      -- CP-element group 73: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/type_cast_1836_konst_delay_trans
      -- CP-element group 73: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/$exit
      -- CP-element group 73: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/$exit
      -- 
    phi_stmt_1832_req_5846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1832_req_5846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(73), ack => phi_stmt_1832_req_0); -- 
    -- Element group convTransposeB_CP_4819_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => convTransposeB_CP_4819_elements(31), ack => convTransposeB_CP_4819_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	31 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1829/SplitProtocol/Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1829/SplitProtocol/Sample/$exit
      -- 
    ra_5863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1829_inst_ack_0, ack => convTransposeB_CP_4819_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	31 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1829/SplitProtocol/Update/ca
      -- CP-element group 75: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1829/SplitProtocol/Update/$exit
      -- 
    ca_5868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1829_inst_ack_1, ack => convTransposeB_CP_4819_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_req
      -- CP-element group 76: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1829/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1829/$exit
      -- CP-element group 76: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/$exit
      -- 
    phi_stmt_1826_req_5869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1826_req_5869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(76), ack => phi_stmt_1826_req_0); -- 
    convTransposeB_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(74) & convTransposeB_CP_4819_elements(75);
      gj_convTransposeB_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	73 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	85 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1684/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(73) & convTransposeB_CP_4819_elements(76);
      gj_convTransposeB_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	70 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/type_cast_1838/SplitProtocol/Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/type_cast_1838/SplitProtocol/Sample/$exit
      -- 
    ra_5889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1838_inst_ack_0, ack => convTransposeB_CP_4819_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	70 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/type_cast_1838/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/type_cast_1838/SplitProtocol/Update/ca
      -- 
    ca_5894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1838_inst_ack_1, ack => convTransposeB_CP_4819_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	84 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/$exit
      -- CP-element group 80: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/type_cast_1838/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_sources/type_cast_1838/$exit
      -- CP-element group 80: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1832/phi_stmt_1832_req
      -- 
    phi_stmt_1832_req_5895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1832_req_5895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(80), ack => phi_stmt_1832_req_1); -- 
    convTransposeB_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(78) & convTransposeB_CP_4819_elements(79);
      gj_convTransposeB_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	70 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1831/SplitProtocol/Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1831/SplitProtocol/Sample/$exit
      -- 
    ra_5912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1831_inst_ack_0, ack => convTransposeB_CP_4819_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	70 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1831/SplitProtocol/Update/ca
      -- CP-element group 82: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1831/SplitProtocol/Update/$exit
      -- 
    ca_5917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1831_inst_ack_1, ack => convTransposeB_CP_4819_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_req
      -- CP-element group 83: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1831/SplitProtocol/$exit
      -- CP-element group 83: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1831/$exit
      -- CP-element group 83: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1826/$exit
      -- 
    phi_stmt_1826_req_5918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1826_req_5918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(83), ack => phi_stmt_1826_req_1); -- 
    convTransposeB_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(81) & convTransposeB_CP_4819_elements(82);
      gj_convTransposeB_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	80 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1684/ifx_xend_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(80) & convTransposeB_CP_4819_elements(83);
      gj_convTransposeB_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  merge  fork  transition  place  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	77 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1684/merge_stmt_1825_PhiReqMerge
      -- CP-element group 85: 	 branch_block_stmt_1684/merge_stmt_1825_PhiAck/$entry
      -- 
    convTransposeB_CP_4819_elements(85) <= OrReduce(convTransposeB_CP_4819_elements(77) & convTransposeB_CP_4819_elements(84));
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1684/merge_stmt_1825_PhiAck/phi_stmt_1826_ack
      -- 
    phi_stmt_1826_ack_5923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1826_ack_0, ack => convTransposeB_CP_4819_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1684/merge_stmt_1825_PhiAck/phi_stmt_1832_ack
      -- 
    phi_stmt_1832_ack_5924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1832_ack_0, ack => convTransposeB_CP_4819_elements(87)); -- 
    -- CP-element group 88:  join  fork  transition  place  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	32 
    -- CP-element group 88: 	33 
    -- CP-element group 88: 	34 
    -- CP-element group 88: 	35 
    -- CP-element group 88:  members (16) 
      -- CP-element group 88: 	 branch_block_stmt_1684/merge_stmt_1825__exit__
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951__entry__
      -- CP-element group 88: 	 branch_block_stmt_1684/merge_stmt_1825_PhiAck/$exit
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/$entry
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1843_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1843_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1843_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1843_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1843_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1843_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1848_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1848_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1848_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1848_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1848_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1684/assign_stmt_1844_to_assign_stmt_1951/type_cast_1848_Update/cr
      -- 
    rr_5436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(88), ack => type_cast_1843_inst_req_0); -- 
    cr_5441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(88), ack => type_cast_1843_inst_req_1); -- 
    rr_5450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(88), ack => type_cast_1848_inst_req_0); -- 
    cr_5455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(88), ack => type_cast_1848_inst_req_1); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(86) & convTransposeB_CP_4819_elements(87);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	59 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Sample/ra
      -- 
    ra_5944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1957_inst_ack_0, ack => convTransposeB_CP_4819_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	59 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Update/ca
      -- CP-element group 90: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Update/$exit
      -- 
    ca_5949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1957_inst_ack_1, ack => convTransposeB_CP_4819_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 91: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/$exit
      -- CP-element group 91: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/$exit
      -- CP-element group 91: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1684/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_req
      -- 
    phi_stmt_1954_req_5950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1954_req_5950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(91), ack => phi_stmt_1954_req_0); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(89) & convTransposeB_CP_4819_elements(90);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  output  delay-element  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	36 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1684/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_req
      -- CP-element group 92: 	 branch_block_stmt_1684/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1960_konst_delay_trans
      -- CP-element group 92: 	 branch_block_stmt_1684/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1684/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1954/$exit
      -- CP-element group 92: 	 branch_block_stmt_1684/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_1954_req_5961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1954_req_5961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(92), ack => phi_stmt_1954_req_1); -- 
    -- Element group convTransposeB_CP_4819_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => convTransposeB_CP_4819_elements(36), ack => convTransposeB_CP_4819_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  merge  transition  place  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1684/merge_stmt_1953_PhiReqMerge
      -- CP-element group 93: 	 branch_block_stmt_1684/merge_stmt_1953_PhiAck/$entry
      -- 
    convTransposeB_CP_4819_elements(93) <= OrReduce(convTransposeB_CP_4819_elements(91) & convTransposeB_CP_4819_elements(92));
    -- CP-element group 94:  fork  transition  place  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	42 
    -- CP-element group 94: 	44 
    -- CP-element group 94: 	46 
    -- CP-element group 94: 	48 
    -- CP-element group 94: 	50 
    -- CP-element group 94: 	52 
    -- CP-element group 94: 	55 
    -- CP-element group 94: 	56 
    -- CP-element group 94: 	57 
    -- CP-element group 94: 	37 
    -- CP-element group 94: 	38 
    -- CP-element group 94: 	40 
    -- CP-element group 94:  members (45) 
      -- CP-element group 94: 	 branch_block_stmt_1684/merge_stmt_1953__exit__
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059__entry__
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_1970_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1684/merge_stmt_1953_PhiAck/phi_stmt_1954_ack
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_1970_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_1970_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_1970_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_1970_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_1970_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1684/merge_stmt_1953_PhiAck/$exit
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2000_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2000_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2000_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2007_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_final_index_sum_regn_update_start
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_final_index_sum_regn_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2006_final_index_sum_regn_Update/req
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2007_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2007_complete/req
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2011_Update/word_access_complete/word_0/cr
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2031_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2031_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2031_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2038_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_final_index_sum_regn_update_start
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_final_index_sum_regn_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/array_obj_ref_2037_final_index_sum_regn_Update/req
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2038_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/addr_of_2038_complete/req
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/ptr_deref_2041_Update/word_access_complete/word_0/cr
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2047_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2047_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2047_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2047_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2047_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1684/assign_stmt_1967_to_assign_stmt_2059/type_cast_2047_Update/cr
      -- 
    phi_stmt_1954_ack_5966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1954_ack_0, ack => convTransposeB_CP_4819_elements(94)); -- 
    rr_5467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(94), ack => type_cast_1970_inst_req_0); -- 
    cr_5472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(94), ack => type_cast_1970_inst_req_1); -- 
    cr_5486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(94), ack => type_cast_2000_inst_req_1); -- 
    req_5517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(94), ack => array_obj_ref_2006_index_offset_req_1); -- 
    req_5532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(94), ack => addr_of_2007_final_reg_req_1); -- 
    cr_5577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(94), ack => ptr_deref_2011_load_0_req_1); -- 
    cr_5596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(94), ack => type_cast_2031_inst_req_1); -- 
    req_5627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(94), ack => array_obj_ref_2037_index_offset_req_1); -- 
    req_5642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(94), ack => addr_of_2038_final_reg_req_1); -- 
    cr_5692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(94), ack => ptr_deref_2041_store_0_req_1); -- 
    rr_5701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(94), ack => type_cast_2047_inst_req_0); -- 
    cr_5706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(94), ack => type_cast_2047_inst_req_1); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	64 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2121/SplitProtocol/Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2121/SplitProtocol/Sample/$exit
      -- 
    ra_6018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2121_inst_ack_0, ack => convTransposeB_CP_4819_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	64 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2121/SplitProtocol/Update/ca
      -- CP-element group 96: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2121/SplitProtocol/Update/$exit
      -- 
    ca_6023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2121_inst_ack_1, ack => convTransposeB_CP_4819_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2121/$exit
      -- CP-element group 97: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2121/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_req
      -- CP-element group 97: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2116/$exit
      -- 
    phi_stmt_2116_req_6024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2116_req_6024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(97), ack => phi_stmt_2116_req_1); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(95) & convTransposeB_CP_4819_elements(96);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	64 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2127/SplitProtocol/Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2127/SplitProtocol/Sample/ra
      -- 
    ra_6041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2127_inst_ack_0, ack => convTransposeB_CP_4819_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	64 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2127/SplitProtocol/Update/ca
      -- CP-element group 99: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2127/SplitProtocol/Update/$exit
      -- 
    ca_6046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2127_inst_ack_1, ack => convTransposeB_CP_4819_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2127/SplitProtocol/$exit
      -- CP-element group 100: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2127/$exit
      -- CP-element group 100: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/$exit
      -- CP-element group 100: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/$exit
      -- CP-element group 100: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_req
      -- 
    phi_stmt_2122_req_6047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2122_req_6047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(100), ack => phi_stmt_2122_req_1); -- 
    convTransposeB_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(98) & convTransposeB_CP_4819_elements(99);
      gj_convTransposeB_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	109 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1684/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(97) & convTransposeB_CP_4819_elements(100);
      gj_convTransposeB_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	66 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2119/SplitProtocol/Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2119/SplitProtocol/Sample/$exit
      -- 
    ra_6067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2119_inst_ack_0, ack => convTransposeB_CP_4819_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	66 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2119/SplitProtocol/Update/ca
      -- CP-element group 103: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2119/SplitProtocol/Update/$exit
      -- 
    ca_6072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2119_inst_ack_1, ack => convTransposeB_CP_4819_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/$exit
      -- CP-element group 104: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2119/$exit
      -- CP-element group 104: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_sources/type_cast_2119/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2116/phi_stmt_2116_req
      -- 
    phi_stmt_2116_req_6073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2116_req_6073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(104), ack => phi_stmt_2116_req_0); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(102) & convTransposeB_CP_4819_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	66 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2125/SplitProtocol/Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2125/SplitProtocol/Sample/$exit
      -- 
    ra_6090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2125_inst_ack_0, ack => convTransposeB_CP_4819_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	66 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2125/SplitProtocol/Update/ca
      -- CP-element group 106: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2125/SplitProtocol/Update/$exit
      -- 
    ca_6095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2125_inst_ack_1, ack => convTransposeB_CP_4819_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_req
      -- CP-element group 107: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2125/$exit
      -- CP-element group 107: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/phi_stmt_2122_sources/type_cast_2125/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2122/$exit
      -- 
    phi_stmt_2122_req_6096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2122_req_6096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(107), ack => phi_stmt_2122_req_0); -- 
    convTransposeB_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(105) & convTransposeB_CP_4819_elements(106);
      gj_convTransposeB_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1684/ifx_xthen79_ifx_xend_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(104) & convTransposeB_CP_4819_elements(107);
      gj_convTransposeB_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  merge  fork  transition  place  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	101 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1684/merge_stmt_2115_PhiReqMerge
      -- CP-element group 109: 	 branch_block_stmt_1684/merge_stmt_2115_PhiAck/$entry
      -- 
    convTransposeB_CP_4819_elements(109) <= OrReduce(convTransposeB_CP_4819_elements(101) & convTransposeB_CP_4819_elements(108));
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1684/merge_stmt_2115_PhiAck/phi_stmt_2116_ack
      -- 
    phi_stmt_2116_ack_6101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2116_ack_0, ack => convTransposeB_CP_4819_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1684/merge_stmt_2115_PhiAck/phi_stmt_2122_ack
      -- 
    phi_stmt_2122_ack_6102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2122_ack_0, ack => convTransposeB_CP_4819_elements(111)); -- 
    -- CP-element group 112:  join  fork  transition  place  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: 	68 
    -- CP-element group 112:  members (10) 
      -- CP-element group 112: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/type_cast_2132_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/type_cast_2132_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/type_cast_2132_Update/cr
      -- CP-element group 112: 	 branch_block_stmt_1684/merge_stmt_2115_PhiAck/$exit
      -- CP-element group 112: 	 branch_block_stmt_1684/merge_stmt_2115__exit__
      -- CP-element group 112: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138__entry__
      -- CP-element group 112: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/type_cast_2132_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/type_cast_2132_update_start_
      -- CP-element group 112: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/type_cast_2132_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1684/assign_stmt_2133_to_assign_stmt_2138/$entry
      -- 
    rr_5793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(112), ack => type_cast_2132_inst_req_0); -- 
    cr_5798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4819_elements(112), ack => type_cast_2132_inst_req_1); -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4819_elements(110) & convTransposeB_CP_4819_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4819_elements(112), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1913_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1934_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1994_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2025_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_1750_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_1750_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom61_2036_resized : std_logic_vector(13 downto 0);
    signal R_idxprom61_2036_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2005_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2005_scaled : std_logic_vector(13 downto 0);
    signal add17_1976 : std_logic_vector(31 downto 0);
    signal add25_1874 : std_logic_vector(31 downto 0);
    signal add36_1889 : std_logic_vector(31 downto 0);
    signal add51_1946 : std_logic_vector(31 downto 0);
    signal add53_1981 : std_logic_vector(31 downto 0);
    signal add66_2054 : std_logic_vector(31 downto 0);
    signal add_1859 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2006_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2006_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2006_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2006_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2006_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2006_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2037_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2037_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2037_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2037_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2037_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2037_root_address : std_logic_vector(13 downto 0);
    signal arrayidx62_2039 : std_logic_vector(31 downto 0);
    signal arrayidx_2008 : std_logic_vector(31 downto 0);
    signal call_1687 : std_logic_vector(15 downto 0);
    signal cmp77_2090 : std_logic_vector(0 downto 0);
    signal cmp89_2138 : std_logic_vector(0 downto 0);
    signal cmp_2059 : std_logic_vector(0 downto 0);
    signal conv12_1844 : std_logic_vector(31 downto 0);
    signal conv15_1849 : std_logic_vector(31 downto 0);
    signal conv22_1736 : std_logic_vector(31 downto 0);
    signal conv27_1755 : std_logic_vector(31 downto 0);
    signal conv33_1769 : std_logic_vector(31 downto 0);
    signal conv46_1915 : std_logic_vector(31 downto 0);
    signal conv49_1936 : std_logic_vector(31 downto 0);
    signal conv65_2048 : std_logic_vector(31 downto 0);
    signal conv75_2085 : std_logic_vector(31 downto 0);
    signal conv84_2113 : std_logic_vector(15 downto 0);
    signal conv86_2133 : std_logic_vector(31 downto 0);
    signal conv9102_1971 : std_logic_vector(31 downto 0);
    signal conv_1710 : std_logic_vector(15 downto 0);
    signal div83_2109 : std_logic_vector(31 downto 0);
    signal div88_1823 : std_logic_vector(31 downto 0);
    signal div_1706 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1813 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1696 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1718 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1728 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1744 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1761 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1777 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1789 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1801 : std_logic_vector(31 downto 0);
    signal idxprom61_2032 : std_logic_vector(63 downto 0);
    signal idxprom_2001 : std_logic_vector(63 downto 0);
    signal inc81_2103 : std_logic_vector(15 downto 0);
    signal inc_2080 : std_logic_vector(15 downto 0);
    signal indvar_1954 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2072 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_2122 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1832 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1826 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2116 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1967 : std_logic_vector(15 downto 0);
    signal mul16_1864 : std_logic_vector(31 downto 0);
    signal mul23_1869 : std_logic_vector(31 downto 0);
    signal mul34_1884 : std_logic_vector(31 downto 0);
    signal mul50_1941 : std_logic_vector(31 downto 0);
    signal mul52_1951 : std_logic_vector(31 downto 0);
    signal mul_1854 : std_logic_vector(31 downto 0);
    signal ptr_deref_1699_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1699_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1699_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1699_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1699_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1721_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1721_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1721_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1721_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1721_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1731_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1731_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1731_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1731_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1731_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1747_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1747_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1747_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1747_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1747_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1764_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1764_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1764_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1764_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1764_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1780_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1780_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1780_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1780_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1780_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1792_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1792_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1792_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1792_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1792_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1804_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1804_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1804_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1804_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1804_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1816_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1816_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1816_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1816_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1816_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2011_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2011_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2011_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2011_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2011_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2041_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2041_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2041_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2041_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2041_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2041_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext103_1927 : std_logic_vector(31 downto 0);
    signal sext105_1987 : std_logic_vector(31 downto 0);
    signal sext106_2018 : std_logic_vector(31 downto 0);
    signal sext_1906 : std_logic_vector(31 downto 0);
    signal shr60_2027 : std_logic_vector(31 downto 0);
    signal shr_1996 : std_logic_vector(31 downto 0);
    signal sub28_1921 : std_logic_vector(31 downto 0);
    signal sub39_1894 : std_logic_vector(31 downto 0);
    signal sub40_1900 : std_logic_vector(31 downto 0);
    signal sub_1879 : std_logic_vector(31 downto 0);
    signal tmp10_1722 : std_logic_vector(31 downto 0);
    signal tmp21_1732 : std_logic_vector(15 downto 0);
    signal tmp24_1748 : std_logic_vector(31 downto 0);
    signal tmp26_1751 : std_logic_vector(15 downto 0);
    signal tmp32_1765 : std_logic_vector(15 downto 0);
    signal tmp35_1781 : std_logic_vector(31 downto 0);
    signal tmp44_1793 : std_logic_vector(31 downto 0);
    signal tmp47_1805 : std_logic_vector(31 downto 0);
    signal tmp57_2012 : std_logic_vector(63 downto 0);
    signal tmp87_1817 : std_logic_vector(31 downto 0);
    signal tmp_1700 : std_logic_vector(31 downto 0);
    signal type_cast_1704_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1821_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1829_wire : std_logic_vector(15 downto 0);
    signal type_cast_1831_wire : std_logic_vector(15 downto 0);
    signal type_cast_1836_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1838_wire : std_logic_vector(15 downto 0);
    signal type_cast_1842_wire : std_logic_vector(31 downto 0);
    signal type_cast_1847_wire : std_logic_vector(31 downto 0);
    signal type_cast_1898_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1904_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1909_wire : std_logic_vector(31 downto 0);
    signal type_cast_1912_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1919_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1925_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1930_wire : std_logic_vector(31 downto 0);
    signal type_cast_1933_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1957_wire : std_logic_vector(15 downto 0);
    signal type_cast_1960_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1965_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1985_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1990_wire : std_logic_vector(31 downto 0);
    signal type_cast_1993_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1999_wire : std_logic_vector(63 downto 0);
    signal type_cast_2016_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2021_wire : std_logic_vector(31 downto 0);
    signal type_cast_2024_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2030_wire : std_logic_vector(63 downto 0);
    signal type_cast_2046_wire : std_logic_vector(31 downto 0);
    signal type_cast_2052_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2070_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2078_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2083_wire : std_logic_vector(31 downto 0);
    signal type_cast_2101_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2107_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2119_wire : std_logic_vector(15 downto 0);
    signal type_cast_2121_wire : std_logic_vector(15 downto 0);
    signal type_cast_2125_wire : std_logic_vector(15 downto 0);
    signal type_cast_2127_wire : std_logic_vector(15 downto 0);
    signal type_cast_2131_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_1750_word_address_0 <= "0";
    array_obj_ref_2006_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2006_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2006_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2006_resized_base_address <= "00000000000000";
    array_obj_ref_2037_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2037_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2037_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2037_resized_base_address <= "00000000000000";
    iNsTr_10_1813 <= "00000000000000000000000000000010";
    iNsTr_2_1696 <= "00000000000000000000000000000011";
    iNsTr_3_1718 <= "00000000000000000000000000000100";
    iNsTr_4_1728 <= "00000000000000000000000000000000";
    iNsTr_5_1744 <= "00000000000000000000000000000011";
    iNsTr_6_1761 <= "00000000000000000000000000000001";
    iNsTr_7_1777 <= "00000000000000000000000000000100";
    iNsTr_8_1789 <= "00000000000000000000000000000100";
    iNsTr_9_1801 <= "00000000000000000000000000000011";
    ptr_deref_1699_word_offset_0 <= "0000000";
    ptr_deref_1721_word_offset_0 <= "0000000";
    ptr_deref_1731_word_offset_0 <= "0";
    ptr_deref_1747_word_offset_0 <= "0000000";
    ptr_deref_1764_word_offset_0 <= "0";
    ptr_deref_1780_word_offset_0 <= "0000000";
    ptr_deref_1792_word_offset_0 <= "0000000";
    ptr_deref_1804_word_offset_0 <= "0000000";
    ptr_deref_1816_word_offset_0 <= "0000000";
    ptr_deref_2011_word_offset_0 <= "00000000000000";
    ptr_deref_2041_word_offset_0 <= "00000000000000";
    type_cast_1704_wire_constant <= "00000000000000000000000000000001";
    type_cast_1821_wire_constant <= "00000000000000000000000000000001";
    type_cast_1836_wire_constant <= "0000000000000000";
    type_cast_1898_wire_constant <= "00000000000000000000000000010000";
    type_cast_1904_wire_constant <= "11111111111111110000000000000000";
    type_cast_1912_wire_constant <= "00000000000000000000000000010000";
    type_cast_1919_wire_constant <= "00000000000000000000000000010000";
    type_cast_1925_wire_constant <= "11111111111111110000000000000000";
    type_cast_1933_wire_constant <= "00000000000000000000000000010000";
    type_cast_1960_wire_constant <= "0000000000000000";
    type_cast_1965_wire_constant <= "0000000000000100";
    type_cast_1985_wire_constant <= "00000000000000000000000000010000";
    type_cast_1993_wire_constant <= "00000000000000000000000000010010";
    type_cast_2016_wire_constant <= "00000000000000000000000000010000";
    type_cast_2024_wire_constant <= "00000000000000000000000000010010";
    type_cast_2052_wire_constant <= "00000000000000000000000000000100";
    type_cast_2070_wire_constant <= "0000000000000001";
    type_cast_2078_wire_constant <= "0000000000000001";
    type_cast_2101_wire_constant <= "0000000000000001";
    type_cast_2107_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_1826: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1829_wire & type_cast_1831_wire;
      req <= phi_stmt_1826_req_0 & phi_stmt_1826_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1826",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1826_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1826,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1826
    phi_stmt_1832: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1836_wire_constant & type_cast_1838_wire;
      req <= phi_stmt_1832_req_0 & phi_stmt_1832_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1832",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1832_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1832,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1832
    phi_stmt_1954: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1957_wire & type_cast_1960_wire_constant;
      req <= phi_stmt_1954_req_0 & phi_stmt_1954_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1954",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1954_ack_0,
          idata => idata,
          odata => indvar_1954,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1954
    phi_stmt_2116: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2119_wire & type_cast_2121_wire;
      req <= phi_stmt_2116_req_0 & phi_stmt_2116_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2116",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2116_ack_0,
          idata => idata,
          odata => input_dim1x_x2_2116,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2116
    phi_stmt_2122: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2125_wire & type_cast_2127_wire;
      req <= phi_stmt_2122_req_0 & phi_stmt_2122_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2122",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2122_ack_0,
          idata => idata,
          odata => input_dim0x_x0_2122,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2122
    addr_of_2007_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2007_final_reg_req_0;
      addr_of_2007_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2007_final_reg_req_1;
      addr_of_2007_final_reg_ack_1<= rack(0);
      addr_of_2007_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2007_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2006_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2008,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2038_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2038_final_reg_req_0;
      addr_of_2038_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2038_final_reg_req_1;
      addr_of_2038_final_reg_ack_1<= rack(0);
      addr_of_2038_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2038_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2037_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx62_2039,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1709_inst_req_0;
      type_cast_1709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1709_inst_req_1;
      type_cast_1709_inst_ack_1<= rack(0);
      type_cast_1709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1706,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1735_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1735_inst_req_0;
      type_cast_1735_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1735_inst_req_1;
      type_cast_1735_inst_ack_1<= rack(0);
      type_cast_1735_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1735_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp21_1732,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_1736,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1754_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1754_inst_req_0;
      type_cast_1754_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1754_inst_req_1;
      type_cast_1754_inst_ack_1<= rack(0);
      type_cast_1754_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1754_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp26_1751,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_1755,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1768_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1768_inst_req_0;
      type_cast_1768_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1768_inst_req_1;
      type_cast_1768_inst_ack_1<= rack(0);
      type_cast_1768_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1768_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp32_1765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_1769,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1829_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1829_inst_req_0;
      type_cast_1829_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1829_inst_req_1;
      type_cast_1829_inst_ack_1<= rack(0);
      type_cast_1829_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1829_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_1710,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1829_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1831_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1831_inst_req_0;
      type_cast_1831_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1831_inst_req_1;
      type_cast_1831_inst_ack_1<= rack(0);
      type_cast_1831_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1831_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2116,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1831_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1838_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1838_inst_req_0;
      type_cast_1838_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1838_inst_req_1;
      type_cast_1838_inst_ack_1<= rack(0);
      type_cast_1838_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1838_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_2122,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1838_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1843_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1843_inst_req_0;
      type_cast_1843_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1843_inst_req_1;
      type_cast_1843_inst_ack_1<= rack(0);
      type_cast_1843_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1843_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1842_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_1844,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1848_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1848_inst_req_0;
      type_cast_1848_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1848_inst_req_1;
      type_cast_1848_inst_ack_1<= rack(0);
      type_cast_1848_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1848_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1847_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_1849,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1909_inst
    process(sext_1906) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_1906(31 downto 0);
      type_cast_1909_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1914_inst
    process(ASHR_i32_i32_1913_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1913_wire(31 downto 0);
      conv46_1915 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1930_inst
    process(sext103_1927) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext103_1927(31 downto 0);
      type_cast_1930_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1935_inst
    process(ASHR_i32_i32_1934_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1934_wire(31 downto 0);
      conv49_1936 <= tmp_var; -- 
    end process;
    type_cast_1957_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1957_inst_req_0;
      type_cast_1957_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1957_inst_req_1;
      type_cast_1957_inst_ack_1<= rack(0);
      type_cast_1957_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1957_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2072,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1957_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1970_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1970_inst_req_0;
      type_cast_1970_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1970_inst_req_1;
      type_cast_1970_inst_ack_1<= rack(0);
      type_cast_1970_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1970_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1967,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9102_1971,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1990_inst
    process(sext105_1987) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext105_1987(31 downto 0);
      type_cast_1990_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1995_inst
    process(ASHR_i32_i32_1994_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1994_wire(31 downto 0);
      shr_1996 <= tmp_var; -- 
    end process;
    type_cast_2000_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2000_inst_req_0;
      type_cast_2000_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2000_inst_req_1;
      type_cast_2000_inst_ack_1<= rack(0);
      type_cast_2000_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2000_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1999_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2001,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2021_inst
    process(sext106_2018) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext106_2018(31 downto 0);
      type_cast_2021_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2026_inst
    process(ASHR_i32_i32_2025_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2025_wire(31 downto 0);
      shr60_2027 <= tmp_var; -- 
    end process;
    type_cast_2031_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2031_inst_req_0;
      type_cast_2031_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2031_inst_req_1;
      type_cast_2031_inst_ack_1<= rack(0);
      type_cast_2031_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2031_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2030_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom61_2032,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2047_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2047_inst_req_0;
      type_cast_2047_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2047_inst_req_1;
      type_cast_2047_inst_ack_1<= rack(0);
      type_cast_2047_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2047_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2046_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2048,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2084_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2084_inst_req_0;
      type_cast_2084_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2084_inst_req_1;
      type_cast_2084_inst_ack_1<= rack(0);
      type_cast_2084_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2084_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2083_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2085,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2112_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2112_inst_req_0;
      type_cast_2112_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2112_inst_req_1;
      type_cast_2112_inst_ack_1<= rack(0);
      type_cast_2112_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2112_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div83_2109,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_2113,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2119_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2119_inst_req_0;
      type_cast_2119_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2119_inst_req_1;
      type_cast_2119_inst_ack_1<= rack(0);
      type_cast_2119_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2119_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv84_2113,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2119_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2121_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2121_inst_req_0;
      type_cast_2121_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2121_inst_req_1;
      type_cast_2121_inst_ack_1<= rack(0);
      type_cast_2121_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2121_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_2080,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2121_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2125_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2125_inst_req_0;
      type_cast_2125_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2125_inst_req_1;
      type_cast_2125_inst_ack_1<= rack(0);
      type_cast_2125_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2125_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc81_2103,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2125_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2127_inst_req_0;
      type_cast_2127_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2127_inst_req_1;
      type_cast_2127_inst_ack_1<= rack(0);
      type_cast_2127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2x_xph_1832,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2127_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2132_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2132_inst_req_0;
      type_cast_2132_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2132_inst_req_1;
      type_cast_2132_inst_ack_1<= rack(0);
      type_cast_2132_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2132_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2131_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_2133,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1750_gather_scatter
    process(LOAD_padding_1750_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1750_data_0;
      ov(15 downto 0) := iv;
      tmp26_1751 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2006_index_1_rename
    process(R_idxprom_2005_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2005_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2005_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2006_index_1_resize
    process(idxprom_2001) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2001;
      ov := iv(13 downto 0);
      R_idxprom_2005_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2006_root_address_inst
    process(array_obj_ref_2006_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2006_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2006_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2037_index_1_rename
    process(R_idxprom61_2036_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom61_2036_resized;
      ov(13 downto 0) := iv;
      R_idxprom61_2036_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2037_index_1_resize
    process(idxprom61_2032) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom61_2032;
      ov := iv(13 downto 0);
      R_idxprom61_2036_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2037_root_address_inst
    process(array_obj_ref_2037_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2037_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2037_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1699_addr_0
    process(ptr_deref_1699_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1699_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1699_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1699_base_resize
    process(iNsTr_2_1696) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1696;
      ov := iv(6 downto 0);
      ptr_deref_1699_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1699_gather_scatter
    process(ptr_deref_1699_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1699_data_0;
      ov(31 downto 0) := iv;
      tmp_1700 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1699_root_address_inst
    process(ptr_deref_1699_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1699_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1699_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1721_addr_0
    process(ptr_deref_1721_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1721_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1721_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1721_base_resize
    process(iNsTr_3_1718) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1718;
      ov := iv(6 downto 0);
      ptr_deref_1721_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1721_gather_scatter
    process(ptr_deref_1721_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1721_data_0;
      ov(31 downto 0) := iv;
      tmp10_1722 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1721_root_address_inst
    process(ptr_deref_1721_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1721_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1721_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1731_addr_0
    process(ptr_deref_1731_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1731_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1731_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1731_base_resize
    process(iNsTr_4_1728) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1728;
      ov := iv(0 downto 0);
      ptr_deref_1731_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1731_gather_scatter
    process(ptr_deref_1731_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1731_data_0;
      ov(15 downto 0) := iv;
      tmp21_1732 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1731_root_address_inst
    process(ptr_deref_1731_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1731_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1731_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1747_addr_0
    process(ptr_deref_1747_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1747_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1747_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1747_base_resize
    process(iNsTr_5_1744) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1744;
      ov := iv(6 downto 0);
      ptr_deref_1747_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1747_gather_scatter
    process(ptr_deref_1747_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1747_data_0;
      ov(31 downto 0) := iv;
      tmp24_1748 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1747_root_address_inst
    process(ptr_deref_1747_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1747_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1747_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1764_addr_0
    process(ptr_deref_1764_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1764_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1764_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1764_base_resize
    process(iNsTr_6_1761) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1761;
      ov := iv(0 downto 0);
      ptr_deref_1764_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1764_gather_scatter
    process(ptr_deref_1764_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1764_data_0;
      ov(15 downto 0) := iv;
      tmp32_1765 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1764_root_address_inst
    process(ptr_deref_1764_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1764_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1764_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1780_addr_0
    process(ptr_deref_1780_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1780_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1780_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1780_base_resize
    process(iNsTr_7_1777) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1777;
      ov := iv(6 downto 0);
      ptr_deref_1780_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1780_gather_scatter
    process(ptr_deref_1780_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1780_data_0;
      ov(31 downto 0) := iv;
      tmp35_1781 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1780_root_address_inst
    process(ptr_deref_1780_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1780_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1780_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1792_addr_0
    process(ptr_deref_1792_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1792_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1792_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1792_base_resize
    process(iNsTr_8_1789) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1789;
      ov := iv(6 downto 0);
      ptr_deref_1792_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1792_gather_scatter
    process(ptr_deref_1792_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1792_data_0;
      ov(31 downto 0) := iv;
      tmp44_1793 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1792_root_address_inst
    process(ptr_deref_1792_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1792_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1792_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1804_addr_0
    process(ptr_deref_1804_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1804_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1804_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1804_base_resize
    process(iNsTr_9_1801) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1801;
      ov := iv(6 downto 0);
      ptr_deref_1804_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1804_gather_scatter
    process(ptr_deref_1804_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1804_data_0;
      ov(31 downto 0) := iv;
      tmp47_1805 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1804_root_address_inst
    process(ptr_deref_1804_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1804_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1804_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1816_addr_0
    process(ptr_deref_1816_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1816_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1816_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1816_base_resize
    process(iNsTr_10_1813) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1813;
      ov := iv(6 downto 0);
      ptr_deref_1816_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1816_gather_scatter
    process(ptr_deref_1816_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1816_data_0;
      ov(31 downto 0) := iv;
      tmp87_1817 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1816_root_address_inst
    process(ptr_deref_1816_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1816_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1816_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2011_addr_0
    process(ptr_deref_2011_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2011_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2011_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2011_base_resize
    process(arrayidx_2008) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2008;
      ov := iv(13 downto 0);
      ptr_deref_2011_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2011_gather_scatter
    process(ptr_deref_2011_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2011_data_0;
      ov(63 downto 0) := iv;
      tmp57_2012 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2011_root_address_inst
    process(ptr_deref_2011_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2011_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2011_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2041_addr_0
    process(ptr_deref_2041_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2041_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2041_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2041_base_resize
    process(arrayidx62_2039) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx62_2039;
      ov := iv(13 downto 0);
      ptr_deref_2041_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2041_gather_scatter
    process(tmp57_2012) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp57_2012;
      ov(63 downto 0) := iv;
      ptr_deref_2041_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2041_root_address_inst
    process(ptr_deref_2041_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2041_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2041_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2060_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2059;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2060_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2060_branch_req_0,
          ack0 => if_stmt_2060_branch_ack_0,
          ack1 => if_stmt_2060_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2091_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_2090;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2091_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2091_branch_req_0,
          ack0 => if_stmt_2091_branch_ack_0,
          ack1 => if_stmt_2091_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2139_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp89_2138;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2139_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2139_branch_req_0,
          ack0 => if_stmt_2139_branch_ack_0,
          ack1 => if_stmt_2139_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2071_inst
    process(indvar_1954) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1954, type_cast_2070_wire_constant, tmp_var);
      indvarx_xnext_2072 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2079_inst
    process(input_dim1x_x1x_xph_1826) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1826, type_cast_2078_wire_constant, tmp_var);
      inc_2080 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2102_inst
    process(input_dim0x_x2x_xph_1832) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_1832, type_cast_2101_wire_constant, tmp_var);
      inc81_2103 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1858_inst
    process(mul_1854, conv12_1844) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_1854, conv12_1844, tmp_var);
      add_1859 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1873_inst
    process(mul23_1869, tmp24_1748) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul23_1869, tmp24_1748, tmp_var);
      add25_1874 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1888_inst
    process(mul34_1884, tmp35_1781) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul34_1884, tmp35_1781, tmp_var);
      add36_1889 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1905_inst
    process(sub40_1900) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub40_1900, type_cast_1904_wire_constant, tmp_var);
      sext_1906 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1926_inst
    process(sub28_1921) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub28_1921, type_cast_1925_wire_constant, tmp_var);
      sext103_1927 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1945_inst
    process(conv46_1915, mul50_1941) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv46_1915, mul50_1941, tmp_var);
      add51_1946 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1975_inst
    process(mul16_1864, conv9102_1971) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul16_1864, conv9102_1971, tmp_var);
      add17_1976 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1980_inst
    process(mul52_1951, conv9102_1971) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul52_1951, conv9102_1971, tmp_var);
      add53_1981 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2053_inst
    process(conv65_2048) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv65_2048, type_cast_2052_wire_constant, tmp_var);
      add66_2054 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1913_inst
    process(type_cast_1909_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1909_wire, type_cast_1912_wire_constant, tmp_var);
      ASHR_i32_i32_1913_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1934_inst
    process(type_cast_1930_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1930_wire, type_cast_1933_wire_constant, tmp_var);
      ASHR_i32_i32_1934_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1994_inst
    process(type_cast_1990_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1990_wire, type_cast_1993_wire_constant, tmp_var);
      ASHR_i32_i32_1994_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2025_inst
    process(type_cast_2021_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2021_wire, type_cast_2024_wire_constant, tmp_var);
      ASHR_i32_i32_2025_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2089_inst
    process(conv75_2085, tmp_1700) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv75_2085, tmp_1700, tmp_var);
      cmp77_2090 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2137_inst
    process(conv86_2133, div88_1823) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv86_2133, div88_1823, tmp_var);
      cmp89_2138 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1705_inst
    process(tmp_1700) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1700, type_cast_1704_wire_constant, tmp_var);
      div_1706 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1822_inst
    process(tmp87_1817) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp87_1817, type_cast_1821_wire_constant, tmp_var);
      div88_1823 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2108_inst
    process(tmp_1700) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1700, type_cast_2107_wire_constant, tmp_var);
      div83_2109 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1966_inst
    process(indvar_1954) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1954, type_cast_1965_wire_constant, tmp_var);
      input_dim2x_x1_1967 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1853_inst
    process(tmp_1700, conv15_1849) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_1700, conv15_1849, tmp_var);
      mul_1854 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1863_inst
    process(add_1859, tmp10_1722) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1859, tmp10_1722, tmp_var);
      mul16_1864 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1868_inst
    process(conv22_1736, conv15_1849) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv22_1736, conv15_1849, tmp_var);
      mul23_1869 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1883_inst
    process(conv33_1769, conv12_1844) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv33_1769, conv12_1844, tmp_var);
      mul34_1884 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1940_inst
    process(tmp47_1805, conv49_1936) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp47_1805, conv49_1936, tmp_var);
      mul50_1941 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1950_inst
    process(add51_1946, tmp44_1793) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add51_1946, tmp44_1793, tmp_var);
      mul52_1951 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1899_inst
    process(sub39_1894) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub39_1894, type_cast_1898_wire_constant, tmp_var);
      sub40_1900 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1920_inst
    process(sub_1879) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_1879, type_cast_1919_wire_constant, tmp_var);
      sub28_1921 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1986_inst
    process(add17_1976) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add17_1976, type_cast_1985_wire_constant, tmp_var);
      sext105_1987 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2017_inst
    process(add53_1981) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add53_1981, type_cast_2016_wire_constant, tmp_var);
      sext106_2018 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1878_inst
    process(add25_1874, conv27_1755) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add25_1874, conv27_1755, tmp_var);
      sub_1879 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1893_inst
    process(add36_1889, conv27_1755) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add36_1889, conv27_1755, tmp_var);
      sub39_1894 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2058_inst
    process(add66_2054, tmp10_1722) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add66_2054, tmp10_1722, tmp_var);
      cmp_2059 <= tmp_var; --
    end process;
    -- shared split operator group (35) : array_obj_ref_2006_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2005_scaled;
      array_obj_ref_2006_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2006_index_offset_req_0;
      array_obj_ref_2006_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2006_index_offset_req_1;
      array_obj_ref_2006_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_2037_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom61_2036_scaled;
      array_obj_ref_2037_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2037_index_offset_req_0;
      array_obj_ref_2037_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2037_index_offset_req_1;
      array_obj_ref_2037_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- unary operator type_cast_1842_inst
    process(input_dim1x_x1x_xph_1826) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_1826, tmp_var);
      type_cast_1842_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1847_inst
    process(input_dim0x_x2x_xph_1832) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_1832, tmp_var);
      type_cast_1847_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1999_inst
    process(shr_1996) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1996, tmp_var);
      type_cast_1999_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2030_inst
    process(shr60_2027) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr60_2027, tmp_var);
      type_cast_2030_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2046_inst
    process(input_dim2x_x1_1967) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_1967, tmp_var);
      type_cast_2046_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2083_inst
    process(inc_2080) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2080, tmp_var);
      type_cast_2083_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2131_inst
    process(input_dim0x_x0_2122) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_2122, tmp_var);
      type_cast_2131_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_1750_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1750_load_0_req_0;
      LOAD_padding_1750_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1750_load_0_req_1;
      LOAD_padding_1750_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1750_word_address_0;
      LOAD_padding_1750_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1699_load_0 ptr_deref_1721_load_0 ptr_deref_1816_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1699_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1721_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1816_load_0_req_0;
      ptr_deref_1699_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1721_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1816_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1699_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1721_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1816_load_0_req_1;
      ptr_deref_1699_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1721_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1816_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1699_word_address_0 & ptr_deref_1721_word_address_0 & ptr_deref_1816_word_address_0;
      ptr_deref_1699_data_0 <= data_out(95 downto 64);
      ptr_deref_1721_data_0 <= data_out(63 downto 32);
      ptr_deref_1816_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1731_load_0 ptr_deref_1764_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1731_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1764_load_0_req_0;
      ptr_deref_1731_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1764_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1731_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1764_load_0_req_1;
      ptr_deref_1731_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1764_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1731_word_address_0 & ptr_deref_1764_word_address_0;
      ptr_deref_1731_data_0 <= data_out(31 downto 16);
      ptr_deref_1764_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1747_load_0 ptr_deref_1780_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1747_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1780_load_0_req_0;
      ptr_deref_1747_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1780_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1747_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1780_load_0_req_1;
      ptr_deref_1747_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1780_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1747_word_address_0 & ptr_deref_1780_word_address_0;
      ptr_deref_1747_data_0 <= data_out(63 downto 32);
      ptr_deref_1780_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1792_load_0 ptr_deref_1804_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1792_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1804_load_0_req_0;
      ptr_deref_1792_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1804_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1792_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1804_load_0_req_1;
      ptr_deref_1792_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1804_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1792_word_address_0 & ptr_deref_1804_word_address_0;
      ptr_deref_1792_data_0 <= data_out(63 downto 32);
      ptr_deref_1804_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2011_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2011_load_0_req_0;
      ptr_deref_2011_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2011_load_0_req_1;
      ptr_deref_2011_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2011_word_address_0;
      ptr_deref_2011_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2041_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2041_store_0_req_0;
      ptr_deref_2041_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2041_store_0_req_1;
      ptr_deref_2041_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2041_word_address_0;
      data_in <= ptr_deref_2041_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1686_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_start_1686_inst_req_0;
      RPIPE_Block1_start_1686_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_start_1686_inst_req_1;
      RPIPE_Block1_start_1686_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1687 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2147_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2147_inst_req_0;
      WPIPE_Block1_done_2147_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2147_inst_req_1;
      WPIPE_Block1_done_2147_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1687;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_6123_start: Boolean;
  signal convTransposeC_CP_6123_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal addr_of_2478_final_reg_ack_0 : boolean;
  signal ptr_deref_2482_load_0_req_1 : boolean;
  signal ptr_deref_2482_load_0_ack_1 : boolean;
  signal type_cast_2441_inst_ack_0 : boolean;
  signal ptr_deref_2275_load_0_req_0 : boolean;
  signal ptr_deref_2275_load_0_ack_1 : boolean;
  signal array_obj_ref_2477_index_offset_req_0 : boolean;
  signal addr_of_2478_final_reg_req_1 : boolean;
  signal type_cast_2502_inst_req_0 : boolean;
  signal addr_of_2478_final_reg_req_0 : boolean;
  signal ptr_deref_2482_load_0_ack_0 : boolean;
  signal type_cast_2314_inst_req_0 : boolean;
  signal type_cast_2314_inst_ack_0 : boolean;
  signal type_cast_2314_inst_req_1 : boolean;
  signal type_cast_2314_inst_ack_1 : boolean;
  signal type_cast_2441_inst_ack_1 : boolean;
  signal type_cast_2319_inst_req_0 : boolean;
  signal type_cast_2319_inst_ack_0 : boolean;
  signal type_cast_2471_inst_req_0 : boolean;
  signal type_cast_2471_inst_ack_0 : boolean;
  signal type_cast_2319_inst_req_1 : boolean;
  signal type_cast_2471_inst_req_1 : boolean;
  signal type_cast_2319_inst_ack_1 : boolean;
  signal array_obj_ref_2477_index_offset_ack_0 : boolean;
  signal type_cast_2502_inst_ack_0 : boolean;
  signal array_obj_ref_2477_index_offset_req_1 : boolean;
  signal addr_of_2478_final_reg_ack_1 : boolean;
  signal array_obj_ref_2477_index_offset_ack_1 : boolean;
  signal type_cast_2502_inst_req_1 : boolean;
  signal type_cast_2502_inst_ack_1 : boolean;
  signal ptr_deref_2287_load_0_req_0 : boolean;
  signal ptr_deref_2287_load_0_ack_0 : boolean;
  signal type_cast_2441_inst_req_1 : boolean;
  signal ptr_deref_2263_load_0_req_1 : boolean;
  signal ptr_deref_2263_load_0_ack_1 : boolean;
  signal ptr_deref_2287_load_0_req_1 : boolean;
  signal ptr_deref_2275_load_0_ack_0 : boolean;
  signal ptr_deref_2287_load_0_ack_1 : boolean;
  signal type_cast_2471_inst_ack_1 : boolean;
  signal ptr_deref_2263_load_0_req_0 : boolean;
  signal type_cast_2441_inst_req_0 : boolean;
  signal ptr_deref_2263_load_0_ack_0 : boolean;
  signal ptr_deref_2275_load_0_req_1 : boolean;
  signal RPIPE_Block2_start_2157_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2157_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2157_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2157_inst_ack_1 : boolean;
  signal ptr_deref_2170_load_0_req_0 : boolean;
  signal ptr_deref_2170_load_0_ack_0 : boolean;
  signal ptr_deref_2170_load_0_req_1 : boolean;
  signal ptr_deref_2170_load_0_ack_1 : boolean;
  signal type_cast_2180_inst_req_0 : boolean;
  signal type_cast_2180_inst_ack_0 : boolean;
  signal type_cast_2180_inst_req_1 : boolean;
  signal type_cast_2180_inst_ack_1 : boolean;
  signal ptr_deref_2192_load_0_req_0 : boolean;
  signal ptr_deref_2192_load_0_ack_0 : boolean;
  signal ptr_deref_2192_load_0_req_1 : boolean;
  signal ptr_deref_2192_load_0_ack_1 : boolean;
  signal ptr_deref_2204_load_0_req_0 : boolean;
  signal ptr_deref_2204_load_0_ack_0 : boolean;
  signal ptr_deref_2204_load_0_req_1 : boolean;
  signal ptr_deref_2204_load_0_ack_1 : boolean;
  signal ptr_deref_2214_load_0_req_0 : boolean;
  signal ptr_deref_2214_load_0_ack_0 : boolean;
  signal ptr_deref_2214_load_0_req_1 : boolean;
  signal ptr_deref_2214_load_0_ack_1 : boolean;
  signal type_cast_2218_inst_req_0 : boolean;
  signal type_cast_2218_inst_ack_0 : boolean;
  signal type_cast_2218_inst_req_1 : boolean;
  signal type_cast_2218_inst_ack_1 : boolean;
  signal ptr_deref_2482_load_0_req_0 : boolean;
  signal ptr_deref_2230_load_0_req_0 : boolean;
  signal ptr_deref_2230_load_0_ack_0 : boolean;
  signal ptr_deref_2230_load_0_req_1 : boolean;
  signal ptr_deref_2230_load_0_ack_1 : boolean;
  signal LOAD_padding_2233_load_0_req_0 : boolean;
  signal LOAD_padding_2233_load_0_ack_0 : boolean;
  signal LOAD_padding_2233_load_0_req_1 : boolean;
  signal LOAD_padding_2233_load_0_ack_1 : boolean;
  signal type_cast_2237_inst_req_0 : boolean;
  signal type_cast_2237_inst_ack_0 : boolean;
  signal type_cast_2237_inst_req_1 : boolean;
  signal type_cast_2237_inst_ack_1 : boolean;
  signal ptr_deref_2247_load_0_req_0 : boolean;
  signal ptr_deref_2247_load_0_ack_0 : boolean;
  signal ptr_deref_2247_load_0_req_1 : boolean;
  signal ptr_deref_2247_load_0_ack_1 : boolean;
  signal type_cast_2251_inst_req_0 : boolean;
  signal type_cast_2251_inst_ack_0 : boolean;
  signal type_cast_2251_inst_req_1 : boolean;
  signal type_cast_2251_inst_ack_1 : boolean;
  signal array_obj_ref_2508_index_offset_req_0 : boolean;
  signal array_obj_ref_2508_index_offset_ack_0 : boolean;
  signal array_obj_ref_2508_index_offset_req_1 : boolean;
  signal array_obj_ref_2508_index_offset_ack_1 : boolean;
  signal addr_of_2509_final_reg_req_0 : boolean;
  signal addr_of_2509_final_reg_ack_0 : boolean;
  signal addr_of_2509_final_reg_req_1 : boolean;
  signal addr_of_2509_final_reg_ack_1 : boolean;
  signal ptr_deref_2512_store_0_req_0 : boolean;
  signal ptr_deref_2512_store_0_ack_0 : boolean;
  signal ptr_deref_2512_store_0_req_1 : boolean;
  signal ptr_deref_2512_store_0_ack_1 : boolean;
  signal type_cast_2518_inst_req_0 : boolean;
  signal type_cast_2518_inst_ack_0 : boolean;
  signal type_cast_2518_inst_req_1 : boolean;
  signal type_cast_2518_inst_ack_1 : boolean;
  signal if_stmt_2531_branch_req_0 : boolean;
  signal if_stmt_2531_branch_ack_1 : boolean;
  signal if_stmt_2531_branch_ack_0 : boolean;
  signal type_cast_2555_inst_req_0 : boolean;
  signal type_cast_2555_inst_ack_0 : boolean;
  signal type_cast_2555_inst_req_1 : boolean;
  signal type_cast_2555_inst_ack_1 : boolean;
  signal type_cast_2564_inst_req_0 : boolean;
  signal type_cast_2564_inst_ack_0 : boolean;
  signal type_cast_2564_inst_req_1 : boolean;
  signal type_cast_2564_inst_ack_1 : boolean;
  signal type_cast_2581_inst_req_0 : boolean;
  signal type_cast_2581_inst_ack_0 : boolean;
  signal type_cast_2581_inst_req_1 : boolean;
  signal type_cast_2581_inst_ack_1 : boolean;
  signal if_stmt_2588_branch_req_0 : boolean;
  signal if_stmt_2588_branch_ack_1 : boolean;
  signal if_stmt_2588_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2596_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2596_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2596_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2596_inst_ack_1 : boolean;
  signal phi_stmt_2297_req_1 : boolean;
  signal type_cast_2309_inst_req_0 : boolean;
  signal type_cast_2309_inst_ack_0 : boolean;
  signal type_cast_2309_inst_req_1 : boolean;
  signal type_cast_2309_inst_ack_1 : boolean;
  signal phi_stmt_2304_req_1 : boolean;
  signal type_cast_2300_inst_req_0 : boolean;
  signal type_cast_2300_inst_ack_0 : boolean;
  signal type_cast_2300_inst_req_1 : boolean;
  signal type_cast_2300_inst_ack_1 : boolean;
  signal phi_stmt_2297_req_0 : boolean;
  signal type_cast_2307_inst_req_0 : boolean;
  signal type_cast_2307_inst_ack_0 : boolean;
  signal type_cast_2307_inst_req_1 : boolean;
  signal type_cast_2307_inst_ack_1 : boolean;
  signal phi_stmt_2304_req_0 : boolean;
  signal phi_stmt_2297_ack_0 : boolean;
  signal phi_stmt_2304_ack_0 : boolean;
  signal type_cast_2431_inst_req_0 : boolean;
  signal type_cast_2431_inst_ack_0 : boolean;
  signal type_cast_2431_inst_req_1 : boolean;
  signal type_cast_2431_inst_ack_1 : boolean;
  signal phi_stmt_2425_req_1 : boolean;
  signal phi_stmt_2425_req_0 : boolean;
  signal phi_stmt_2425_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_6123_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_6123_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_6123_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_6123_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_6123: Block -- control-path 
    signal convTransposeC_CP_6123_elements: BooleanArray(92 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_6123_elements(0) <= convTransposeC_CP_6123_start;
    convTransposeC_CP_6123_symbol <= convTransposeC_CP_6123_elements(70);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2155/$entry
      -- CP-element group 0: 	 branch_block_stmt_2155/branch_block_stmt_2155__entry__
      -- CP-element group 0: 	 branch_block_stmt_2155/assign_stmt_2158__entry__
      -- CP-element group 0: 	 branch_block_stmt_2155/assign_stmt_2158/$entry
      -- CP-element group 0: 	 branch_block_stmt_2155/assign_stmt_2158/RPIPE_Block2_start_2157_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2155/assign_stmt_2158/RPIPE_Block2_start_2157_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2155/assign_stmt_2158/RPIPE_Block2_start_2157_Sample/rr
      -- 
    rr_6171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(0), ack => RPIPE_Block2_start_2157_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2155/assign_stmt_2158/RPIPE_Block2_start_2157_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2155/assign_stmt_2158/RPIPE_Block2_start_2157_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2155/assign_stmt_2158/RPIPE_Block2_start_2157_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2155/assign_stmt_2158/RPIPE_Block2_start_2157_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2155/assign_stmt_2158/RPIPE_Block2_start_2157_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2155/assign_stmt_2158/RPIPE_Block2_start_2157_Update/cr
      -- 
    ra_6172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2157_inst_ack_0, ack => convTransposeC_CP_6123_elements(1)); -- 
    cr_6176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(1), ack => RPIPE_Block2_start_2157_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (265) 
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2158__exit__
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294__entry__
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2158/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2158/RPIPE_Block2_start_2157_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2158/RPIPE_Block2_start_2157_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2158/RPIPE_Block2_start_2157_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2180_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2180_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2180_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2218_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2218_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2218_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2237_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2237_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2237_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2251_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2251_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2251_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_sample_start_
      -- 
    ca_6177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2157_inst_ack_1, ack => convTransposeC_CP_6123_elements(2)); -- 
    rr_6652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2275_load_0_req_0); -- 
    rr_6702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2287_load_0_req_0); -- 
    cr_6613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2263_load_0_req_1); -- 
    cr_6713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2287_load_0_req_1); -- 
    rr_6602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2263_load_0_req_0); -- 
    cr_6663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2275_load_0_req_1); -- 
    rr_6213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2170_load_0_req_0); -- 
    cr_6224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2170_load_0_req_1); -- 
    cr_6243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => type_cast_2180_inst_req_1); -- 
    rr_6277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2192_load_0_req_0); -- 
    cr_6288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2192_load_0_req_1); -- 
    rr_6327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2204_load_0_req_0); -- 
    cr_6338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2204_load_0_req_1); -- 
    rr_6377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2214_load_0_req_0); -- 
    cr_6388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2214_load_0_req_1); -- 
    cr_6407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => type_cast_2218_inst_req_1); -- 
    rr_6441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2230_load_0_req_0); -- 
    cr_6452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2230_load_0_req_1); -- 
    rr_6474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => LOAD_padding_2233_load_0_req_0); -- 
    cr_6485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => LOAD_padding_2233_load_0_req_1); -- 
    cr_6504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => type_cast_2237_inst_req_1); -- 
    rr_6538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2247_load_0_req_0); -- 
    cr_6549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => ptr_deref_2247_load_0_req_1); -- 
    cr_6568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(2), ack => type_cast_2251_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Sample/word_access_start/word_0/ra
      -- 
    ra_6214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2170_load_0_ack_0, ack => convTransposeC_CP_6123_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Update/ptr_deref_2170_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Update/ptr_deref_2170_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Update/ptr_deref_2170_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2170_Update/ptr_deref_2170_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2180_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2180_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2180_Sample/rr
      -- 
    ca_6225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2170_load_0_ack_1, ack => convTransposeC_CP_6123_elements(4)); -- 
    rr_6238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(4), ack => type_cast_2180_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2180_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2180_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2180_Sample/ra
      -- 
    ra_6239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2180_inst_ack_0, ack => convTransposeC_CP_6123_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	31 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2180_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2180_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2180_Update/ca
      -- 
    ca_6244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2180_inst_ack_1, ack => convTransposeC_CP_6123_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Sample/word_access_start/word_0/ra
      -- 
    ra_6278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2192_load_0_ack_0, ack => convTransposeC_CP_6123_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	31 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Update/ptr_deref_2192_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Update/ptr_deref_2192_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Update/ptr_deref_2192_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2192_Update/ptr_deref_2192_Merge/merge_ack
      -- 
    ca_6289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2192_load_0_ack_1, ack => convTransposeC_CP_6123_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Sample/word_access_start/word_0/ra
      -- 
    ra_6328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2204_load_0_ack_0, ack => convTransposeC_CP_6123_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	31 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Update/ptr_deref_2204_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Update/ptr_deref_2204_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Update/ptr_deref_2204_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2204_Update/ptr_deref_2204_Merge/merge_ack
      -- 
    ca_6339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2204_load_0_ack_1, ack => convTransposeC_CP_6123_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Sample/word_access_start/word_0/ra
      -- 
    ra_6378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2214_load_0_ack_0, ack => convTransposeC_CP_6123_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (12) 
      -- CP-element group 12: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Update/ptr_deref_2214_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Update/ptr_deref_2214_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Update/ptr_deref_2214_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2214_Update/ptr_deref_2214_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2218_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2218_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2218_Sample/rr
      -- 
    ca_6389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2214_load_0_ack_1, ack => convTransposeC_CP_6123_elements(12)); -- 
    rr_6402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(12), ack => type_cast_2218_inst_req_0); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2218_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2218_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2218_Sample/ra
      -- 
    ra_6403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2218_inst_ack_0, ack => convTransposeC_CP_6123_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	31 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2218_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2218_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2218_Update/ca
      -- 
    ca_6408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2218_inst_ack_1, ack => convTransposeC_CP_6123_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Sample/word_access_start/word_0/ra
      -- 
    ra_6442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2230_load_0_ack_0, ack => convTransposeC_CP_6123_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	31 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Update/ptr_deref_2230_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Update/ptr_deref_2230_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Update/ptr_deref_2230_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2230_Update/ptr_deref_2230_Merge/merge_ack
      -- 
    ca_6453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2230_load_0_ack_1, ack => convTransposeC_CP_6123_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Sample/word_access_start/word_0/ra
      -- 
    ra_6475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2233_load_0_ack_0, ack => convTransposeC_CP_6123_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (12) 
      -- CP-element group 18: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Update/LOAD_padding_2233_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Update/LOAD_padding_2233_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Update/LOAD_padding_2233_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/LOAD_padding_2233_Update/LOAD_padding_2233_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2237_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2237_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2237_Sample/rr
      -- 
    ca_6486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2233_load_0_ack_1, ack => convTransposeC_CP_6123_elements(18)); -- 
    rr_6499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(18), ack => type_cast_2237_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2237_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2237_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2237_Sample/ra
      -- 
    ra_6500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2237_inst_ack_0, ack => convTransposeC_CP_6123_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	31 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2237_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2237_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2237_Update/ca
      -- 
    ca_6505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2237_inst_ack_1, ack => convTransposeC_CP_6123_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Sample/word_access_start/word_0/ra
      -- 
    ra_6539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2247_load_0_ack_0, ack => convTransposeC_CP_6123_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (12) 
      -- CP-element group 22: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Update/ptr_deref_2247_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Update/ptr_deref_2247_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Update/ptr_deref_2247_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2247_Update/ptr_deref_2247_Merge/merge_ack
      -- CP-element group 22: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2251_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2251_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2251_Sample/rr
      -- 
    ca_6550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2247_load_0_ack_1, ack => convTransposeC_CP_6123_elements(22)); -- 
    rr_6563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(22), ack => type_cast_2251_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2251_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2251_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2251_Sample/ra
      -- 
    ra_6564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2251_inst_ack_0, ack => convTransposeC_CP_6123_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	31 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2251_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2251_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/type_cast_2251_Update/ca
      -- 
    ca_6569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2251_inst_ack_1, ack => convTransposeC_CP_6123_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Sample/word_access_start/word_0/ra
      -- CP-element group 25: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_sample_completed_
      -- 
    ra_6603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2263_load_0_ack_0, ack => convTransposeC_CP_6123_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Update/ptr_deref_2263_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Update/ptr_deref_2263_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Update/ptr_deref_2263_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Update/ptr_deref_2263_Merge/merge_ack
      -- CP-element group 26: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2263_update_completed_
      -- 
    ca_6614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2263_load_0_ack_1, ack => convTransposeC_CP_6123_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Sample/word_access_start/word_0/ra
      -- CP-element group 27: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Sample/word_access_start/$exit
      -- 
    ra_6653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2275_load_0_ack_0, ack => convTransposeC_CP_6123_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Update/ptr_deref_2275_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Update/ptr_deref_2275_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Update/ptr_deref_2275_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Update/ptr_deref_2275_Merge/merge_ack
      -- CP-element group 28: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2275_Update/word_access_complete/word_0/$exit
      -- 
    ca_6664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2275_load_0_ack_1, ack => convTransposeC_CP_6123_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Sample/word_access_start/word_0/ra
      -- CP-element group 29: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Sample/word_access_start/$exit
      -- 
    ra_6703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2287_load_0_ack_0, ack => convTransposeC_CP_6123_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Update/ptr_deref_2287_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Update/ptr_deref_2287_Merge/$exit
      -- CP-element group 30: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Update/ptr_deref_2287_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Update/ptr_deref_2287_Merge/merge_ack
      -- CP-element group 30: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/ptr_deref_2287_update_completed_
      -- 
    ca_6714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2287_load_0_ack_1, ack => convTransposeC_CP_6123_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	10 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	16 
    -- CP-element group 31: 	14 
    -- CP-element group 31: 	24 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	20 
    -- CP-element group 31: 	6 
    -- CP-element group 31: 	8 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	73 
    -- CP-element group 31: 	71 
    -- CP-element group 31: 	72 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294__exit__
      -- CP-element group 31: 	 branch_block_stmt_2155/assign_stmt_2167_to_assign_stmt_2294/$exit
      -- CP-element group 31: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/$entry
      -- CP-element group 31: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/$entry
      -- CP-element group 31: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/$entry
      -- CP-element group 31: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/cr
      -- 
    rr_7131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(31), ack => type_cast_2309_inst_req_0); -- 
    cr_7136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(31), ack => type_cast_2309_inst_req_1); -- 
    convTransposeC_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeC_CP_6123_elements(10) & convTransposeC_CP_6123_elements(30) & convTransposeC_CP_6123_elements(16) & convTransposeC_CP_6123_elements(14) & convTransposeC_CP_6123_elements(24) & convTransposeC_CP_6123_elements(28) & convTransposeC_CP_6123_elements(26) & convTransposeC_CP_6123_elements(20) & convTransposeC_CP_6123_elements(6) & convTransposeC_CP_6123_elements(8);
      gj_convTransposeC_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6123_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	86 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2314_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2314_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2314_sample_completed_
      -- 
    ra_6731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2314_inst_ack_0, ack => convTransposeC_CP_6123_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	86 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2314_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2314_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2314_Update/ca
      -- 
    ca_6736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2314_inst_ack_1, ack => convTransposeC_CP_6123_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	86 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2319_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2319_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2319_Sample/ra
      -- 
    ra_6745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2319_inst_ack_0, ack => convTransposeC_CP_6123_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	86 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2319_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2319_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2319_Update/ca
      -- 
    ca_6750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2319_inst_ack_1, ack => convTransposeC_CP_6123_elements(35)); -- 
    -- CP-element group 36:  join  transition  place  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	33 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	90 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_2155/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 36: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422__exit__
      -- CP-element group 36: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/$exit
      -- CP-element group 36: 	 branch_block_stmt_2155/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_2155/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2425/$entry
      -- CP-element group 36: 	 branch_block_stmt_2155/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/$entry
      -- 
    convTransposeC_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6123_elements(33) & convTransposeC_CP_6123_elements(35);
      gj_convTransposeC_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6123_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	92 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2441_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2441_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2441_Sample/$exit
      -- 
    ra_6762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2441_inst_ack_0, ack => convTransposeC_CP_6123_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	92 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	47 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2502_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2502_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2441_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2471_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2471_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2471_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2441_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2502_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2441_Update/$exit
      -- 
    ca_6767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2441_inst_ack_1, ack => convTransposeC_CP_6123_elements(38)); -- 
    rr_6775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(38), ack => type_cast_2471_inst_req_0); -- 
    rr_6885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(38), ack => type_cast_2502_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2471_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2471_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2471_Sample/ra
      -- 
    ra_6776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2471_inst_ack_0, ack => convTransposeC_CP_6123_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	92 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (16) 
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_index_scale_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_index_scale_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_index_scale_1/scale_rename_req
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_final_index_sum_regn_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_final_index_sum_regn_Sample/req
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_index_computed_1
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2471_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2471_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_index_resize_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_index_resize_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_index_scale_1/scale_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_index_resize_1/index_resize_req
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_index_resized_1
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2471_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_index_scaled_1
      -- CP-element group 40: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_index_resize_1/index_resize_ack
      -- 
    ca_6781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2471_inst_ack_1, ack => convTransposeC_CP_6123_elements(40)); -- 
    req_6806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(40), ack => array_obj_ref_2477_index_offset_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_final_index_sum_regn_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_final_index_sum_regn_Sample/ack
      -- CP-element group 41: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_final_index_sum_regn_sample_complete
      -- 
    ack_6807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2477_index_offset_ack_0, ack => convTransposeC_CP_6123_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	92 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (11) 
      -- CP-element group 42: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_offset_calculated
      -- CP-element group 42: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2478_request/req
      -- CP-element group 42: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_final_index_sum_regn_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_final_index_sum_regn_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2478_request/$entry
      -- CP-element group 42: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2478_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_root_address_calculated
      -- 
    ack_6812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2477_index_offset_ack_1, ack => convTransposeC_CP_6123_elements(42)); -- 
    req_6821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(42), ack => addr_of_2478_final_reg_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2478_request/ack
      -- CP-element group 43: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2478_request/$exit
      -- CP-element group 43: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2478_sample_completed_
      -- 
    ack_6822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2478_final_reg_ack_0, ack => convTransposeC_CP_6123_elements(43)); -- 
    -- CP-element group 44:  join  fork  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	92 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (24) 
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_base_addr_resize/base_resize_req
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2478_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_word_addrgen/$entry
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_word_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2478_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_word_addrgen/$exit
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_word_addrgen/root_register_req
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_word_addrgen/root_register_ack
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2478_complete/ack
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Sample/word_access_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_base_address_resized
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_base_addr_resize/base_resize_ack
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_base_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_base_addr_resize/$entry
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_base_addr_resize/$exit
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Sample/word_access_start/word_0/rr
      -- 
    ack_6827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2478_final_reg_ack_1, ack => convTransposeC_CP_6123_elements(44)); -- 
    rr_6860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(44), ack => ptr_deref_2482_load_0_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Sample/word_access_start/word_0/ra
      -- CP-element group 45: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Sample/word_access_start/word_0/$exit
      -- 
    ra_6861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2482_load_0_ack_0, ack => convTransposeC_CP_6123_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	92 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	53 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Update/word_access_complete/word_0/ca
      -- CP-element group 46: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Update/ptr_deref_2482_Merge/$entry
      -- CP-element group 46: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Update/ptr_deref_2482_Merge/$exit
      -- CP-element group 46: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Update/ptr_deref_2482_Merge/merge_req
      -- CP-element group 46: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Update/ptr_deref_2482_Merge/merge_ack
      -- CP-element group 46: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_update_completed_
      -- 
    ca_6872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2482_load_0_ack_1, ack => convTransposeC_CP_6123_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	38 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2502_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2502_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2502_Sample/ra
      -- 
    ra_6886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2502_inst_ack_0, ack => convTransposeC_CP_6123_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	92 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (16) 
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2502_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2502_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2502_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_index_resized_1
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_index_scaled_1
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_index_computed_1
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_index_resize_1/index_resize_req
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_index_resize_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_index_resize_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_index_resize_1/index_resize_ack
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_index_scale_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_index_scale_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_index_scale_1/scale_rename_req
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_index_scale_1/scale_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_final_index_sum_regn_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_final_index_sum_regn_Sample/req
      -- 
    ca_6891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2502_inst_ack_1, ack => convTransposeC_CP_6123_elements(48)); -- 
    req_6916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(48), ack => array_obj_ref_2508_index_offset_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_final_index_sum_regn_sample_complete
      -- CP-element group 49: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_final_index_sum_regn_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_final_index_sum_regn_Sample/ack
      -- 
    ack_6917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2508_index_offset_ack_0, ack => convTransposeC_CP_6123_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	92 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (11) 
      -- CP-element group 50: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2509_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_offset_calculated
      -- CP-element group 50: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2509_request/$entry
      -- CP-element group 50: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_final_index_sum_regn_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_final_index_sum_regn_Update/ack
      -- CP-element group 50: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2509_request/req
      -- 
    ack_6922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2508_index_offset_ack_1, ack => convTransposeC_CP_6123_elements(50)); -- 
    req_6931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(50), ack => addr_of_2509_final_reg_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2509_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2509_request/$exit
      -- CP-element group 51: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2509_request/ack
      -- 
    ack_6932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2509_final_reg_ack_0, ack => convTransposeC_CP_6123_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	92 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (19) 
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2509_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2509_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2509_complete/ack
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_word_addrgen/root_register_ack
      -- 
    ack_6937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2509_final_reg_ack_1, ack => convTransposeC_CP_6123_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	46 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Sample/ptr_deref_2512_Split/$entry
      -- CP-element group 53: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Sample/ptr_deref_2512_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Sample/ptr_deref_2512_Split/split_req
      -- CP-element group 53: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Sample/ptr_deref_2512_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Sample/word_access_start/word_0/rr
      -- 
    rr_6975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(53), ack => ptr_deref_2512_store_0_req_0); -- 
    convTransposeC_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6123_elements(46) & convTransposeC_CP_6123_elements(52);
      gj_convTransposeC_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6123_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Sample/word_access_start/word_0/ra
      -- 
    ra_6976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2512_store_0_ack_0, ack => convTransposeC_CP_6123_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	92 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Update/word_access_complete/word_0/ca
      -- 
    ca_6987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2512_store_0_ack_1, ack => convTransposeC_CP_6123_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	92 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2518_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2518_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2518_Sample/ra
      -- 
    ra_6996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2518_inst_ack_0, ack => convTransposeC_CP_6123_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	92 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2518_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2518_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2518_Update/ca
      -- 
    ca_7001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2518_inst_ack_1, ack => convTransposeC_CP_6123_elements(57)); -- 
    -- CP-element group 58:  branch  join  transition  place  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	55 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (10) 
      -- CP-element group 58: 	 branch_block_stmt_2155/R_cmp_2532_place
      -- CP-element group 58: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530__exit__
      -- CP-element group 58: 	 branch_block_stmt_2155/if_stmt_2531__entry__
      -- CP-element group 58: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/$exit
      -- CP-element group 58: 	 branch_block_stmt_2155/if_stmt_2531_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2155/if_stmt_2531_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_2155/if_stmt_2531_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_2155/if_stmt_2531_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_2155/if_stmt_2531_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2155/if_stmt_2531_else_link/$entry
      -- 
    branch_req_7009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(58), ack => if_stmt_2531_branch_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_6123_elements(41) & convTransposeC_CP_6123_elements(55) & convTransposeC_CP_6123_elements(57) & convTransposeC_CP_6123_elements(49);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6123_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	87 
    -- CP-element group 59: 	88 
    -- CP-element group 59:  members (24) 
      -- CP-element group 59: 	 branch_block_stmt_2155/whilex_xbody_ifx_xthen
      -- CP-element group 59: 	 branch_block_stmt_2155/assign_stmt_2543__exit__
      -- CP-element group 59: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody
      -- CP-element group 59: 	 branch_block_stmt_2155/merge_stmt_2537__exit__
      -- CP-element group 59: 	 branch_block_stmt_2155/assign_stmt_2543__entry__
      -- CP-element group 59: 	 branch_block_stmt_2155/if_stmt_2531_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_2155/if_stmt_2531_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_2155/assign_stmt_2543/$entry
      -- CP-element group 59: 	 branch_block_stmt_2155/assign_stmt_2543/$exit
      -- CP-element group 59: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/$entry
      -- CP-element group 59: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/$entry
      -- CP-element group 59: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Update/cr
      -- CP-element group 59: 	 branch_block_stmt_2155/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_2155/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_2155/merge_stmt_2537_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_2155/merge_stmt_2537_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_2155/merge_stmt_2537_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_2155/merge_stmt_2537_PhiAck/dummy
      -- 
    if_choice_transition_7014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2531_branch_ack_1, ack => convTransposeC_CP_6123_elements(59)); -- 
    rr_7212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(59), ack => type_cast_2431_inst_req_0); -- 
    cr_7217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(59), ack => type_cast_2431_inst_req_1); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	66 
    -- CP-element group 60: 	64 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (24) 
      -- CP-element group 60: 	 branch_block_stmt_2155/whilex_xbody_ifx_xelse
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587__entry__
      -- CP-element group 60: 	 branch_block_stmt_2155/merge_stmt_2545__exit__
      -- CP-element group 60: 	 branch_block_stmt_2155/if_stmt_2531_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_2155/if_stmt_2531_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/$entry
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2555_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2555_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2555_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2555_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2555_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2555_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2564_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2564_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2564_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2581_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2581_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2581_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2155/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_2155/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_2155/merge_stmt_2545_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_2155/merge_stmt_2545_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_2155/merge_stmt_2545_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_2155/merge_stmt_2545_PhiAck/dummy
      -- 
    else_choice_transition_7018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2531_branch_ack_0, ack => convTransposeC_CP_6123_elements(60)); -- 
    rr_7034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(60), ack => type_cast_2555_inst_req_0); -- 
    cr_7039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(60), ack => type_cast_2555_inst_req_1); -- 
    cr_7053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(60), ack => type_cast_2564_inst_req_1); -- 
    cr_7067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(60), ack => type_cast_2581_inst_req_1); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2555_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2555_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2555_Sample/ra
      -- 
    ra_7035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2555_inst_ack_0, ack => convTransposeC_CP_6123_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2555_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2555_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2555_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2564_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2564_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2564_Sample/rr
      -- 
    ca_7040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2555_inst_ack_1, ack => convTransposeC_CP_6123_elements(62)); -- 
    rr_7048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(62), ack => type_cast_2564_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2564_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2564_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2564_Sample/ra
      -- 
    ra_7049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2564_inst_ack_0, ack => convTransposeC_CP_6123_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	60 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2564_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2564_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2564_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2581_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2581_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2581_Sample/rr
      -- 
    ca_7054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2564_inst_ack_1, ack => convTransposeC_CP_6123_elements(64)); -- 
    rr_7062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(64), ack => type_cast_2581_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2581_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2581_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2581_Sample/ra
      -- 
    ra_7063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2581_inst_ack_0, ack => convTransposeC_CP_6123_elements(65)); -- 
    -- CP-element group 66:  branch  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	60 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (13) 
      -- CP-element group 66: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587__exit__
      -- CP-element group 66: 	 branch_block_stmt_2155/if_stmt_2588__entry__
      -- CP-element group 66: 	 branch_block_stmt_2155/R_cmp87_2589_place
      -- CP-element group 66: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/$exit
      -- CP-element group 66: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2581_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2581_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2155/assign_stmt_2551_to_assign_stmt_2587/type_cast_2581_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_2155/if_stmt_2588_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2155/if_stmt_2588_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2155/if_stmt_2588_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2155/if_stmt_2588_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2155/if_stmt_2588_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2155/if_stmt_2588_else_link/$entry
      -- 
    ca_7068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2581_inst_ack_1, ack => convTransposeC_CP_6123_elements(66)); -- 
    branch_req_7076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(66), ack => if_stmt_2588_branch_req_0); -- 
    -- CP-element group 67:  merge  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (15) 
      -- CP-element group 67: 	 branch_block_stmt_2155/merge_stmt_2594__exit__
      -- CP-element group 67: 	 branch_block_stmt_2155/assign_stmt_2598__entry__
      -- CP-element group 67: 	 branch_block_stmt_2155/if_stmt_2588_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2155/if_stmt_2588_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2155/ifx_xelse_whilex_xend
      -- CP-element group 67: 	 branch_block_stmt_2155/assign_stmt_2598/$entry
      -- CP-element group 67: 	 branch_block_stmt_2155/assign_stmt_2598/WPIPE_Block2_done_2596_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_2155/assign_stmt_2598/WPIPE_Block2_done_2596_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2155/assign_stmt_2598/WPIPE_Block2_done_2596_Sample/req
      -- CP-element group 67: 	 branch_block_stmt_2155/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2155/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2155/merge_stmt_2594_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2155/merge_stmt_2594_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2155/merge_stmt_2594_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2155/merge_stmt_2594_PhiAck/dummy
      -- 
    if_choice_transition_7081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2588_branch_ack_1, ack => convTransposeC_CP_6123_elements(67)); -- 
    req_7098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(67), ack => WPIPE_Block2_done_2596_inst_req_0); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	76 
    -- CP-element group 68: 	77 
    -- CP-element group 68: 	79 
    -- CP-element group 68: 	80 
    -- CP-element group 68:  members (20) 
      -- CP-element group 68: 	 branch_block_stmt_2155/if_stmt_2588_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_2155/if_stmt_2588_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/$entry
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/$entry
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/$entry
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/$entry
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2588_branch_ack_0, ack => convTransposeC_CP_6123_elements(68)); -- 
    rr_7157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(68), ack => type_cast_2300_inst_req_0); -- 
    cr_7162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(68), ack => type_cast_2300_inst_req_1); -- 
    rr_7180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(68), ack => type_cast_2307_inst_req_0); -- 
    cr_7185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(68), ack => type_cast_2307_inst_req_1); -- 
    -- CP-element group 69:  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_2155/assign_stmt_2598/WPIPE_Block2_done_2596_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2155/assign_stmt_2598/WPIPE_Block2_done_2596_update_start_
      -- CP-element group 69: 	 branch_block_stmt_2155/assign_stmt_2598/WPIPE_Block2_done_2596_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2155/assign_stmt_2598/WPIPE_Block2_done_2596_Sample/ack
      -- CP-element group 69: 	 branch_block_stmt_2155/assign_stmt_2598/WPIPE_Block2_done_2596_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2155/assign_stmt_2598/WPIPE_Block2_done_2596_Update/req
      -- 
    ack_7099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2596_inst_ack_0, ack => convTransposeC_CP_6123_elements(69)); -- 
    req_7103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(69), ack => WPIPE_Block2_done_2596_inst_req_1); -- 
    -- CP-element group 70:  transition  place  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (16) 
      -- CP-element group 70: 	 $exit
      -- CP-element group 70: 	 branch_block_stmt_2155/$exit
      -- CP-element group 70: 	 branch_block_stmt_2155/branch_block_stmt_2155__exit__
      -- CP-element group 70: 	 branch_block_stmt_2155/assign_stmt_2598__exit__
      -- CP-element group 70: 	 branch_block_stmt_2155/return__
      -- CP-element group 70: 	 branch_block_stmt_2155/merge_stmt_2600__exit__
      -- CP-element group 70: 	 branch_block_stmt_2155/assign_stmt_2598/$exit
      -- CP-element group 70: 	 branch_block_stmt_2155/assign_stmt_2598/WPIPE_Block2_done_2596_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2155/assign_stmt_2598/WPIPE_Block2_done_2596_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2155/assign_stmt_2598/WPIPE_Block2_done_2596_Update/ack
      -- CP-element group 70: 	 branch_block_stmt_2155/return___PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_2155/return___PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2155/merge_stmt_2600_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2155/merge_stmt_2600_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2155/merge_stmt_2600_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2155/merge_stmt_2600_PhiAck/dummy
      -- 
    ack_7104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2596_inst_ack_1, ack => convTransposeC_CP_6123_elements(70)); -- 
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	75 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/$exit
      -- CP-element group 71: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2303_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_req
      -- 
    phi_stmt_2297_req_7115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2297_req_7115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(71), ack => phi_stmt_2297_req_1); -- 
    -- Element group convTransposeC_CP_6123_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => convTransposeC_CP_6123_elements(31), ack => convTransposeC_CP_6123_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	31 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Sample/ra
      -- 
    ra_7132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2309_inst_ack_0, ack => convTransposeC_CP_6123_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	31 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/Update/ca
      -- 
    ca_7137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2309_inst_ack_1, ack => convTransposeC_CP_6123_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/$exit
      -- CP-element group 74: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/$exit
      -- CP-element group 74: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2309/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_req
      -- 
    phi_stmt_2304_req_7138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2304_req_7138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(74), ack => phi_stmt_2304_req_1); -- 
    convTransposeC_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6123_elements(73) & convTransposeC_CP_6123_elements(72);
      gj_convTransposeC_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6123_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: 	71 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	83 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_2155/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6123_elements(74) & convTransposeC_CP_6123_elements(71);
      gj_convTransposeC_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6123_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	68 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Sample/ra
      -- 
    ra_7158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2300_inst_ack_0, ack => convTransposeC_CP_6123_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	68 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Update/ca
      -- 
    ca_7163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2300_inst_ack_1, ack => convTransposeC_CP_6123_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	82 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/$exit
      -- CP-element group 78: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/$exit
      -- CP-element group 78: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/$exit
      -- CP-element group 78: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2297/phi_stmt_2297_req
      -- 
    phi_stmt_2297_req_7164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2297_req_7164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(78), ack => phi_stmt_2297_req_0); -- 
    convTransposeC_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6123_elements(76) & convTransposeC_CP_6123_elements(77);
      gj_convTransposeC_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6123_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	68 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Sample/ra
      -- 
    ra_7181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2307_inst_ack_0, ack => convTransposeC_CP_6123_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	68 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/Update/ca
      -- 
    ca_7186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2307_inst_ack_1, ack => convTransposeC_CP_6123_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/$exit
      -- CP-element group 81: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/$exit
      -- CP-element group 81: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_sources/type_cast_2307/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2304/phi_stmt_2304_req
      -- 
    phi_stmt_2304_req_7187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2304_req_7187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(81), ack => phi_stmt_2304_req_0); -- 
    convTransposeC_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6123_elements(79) & convTransposeC_CP_6123_elements(80);
      gj_convTransposeC_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6123_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  transition  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_2155/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6123_elements(78) & convTransposeC_CP_6123_elements(81);
      gj_convTransposeC_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6123_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  merge  fork  transition  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	75 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2155/merge_stmt_2296_PhiReqMerge
      -- CP-element group 83: 	 branch_block_stmt_2155/merge_stmt_2296_PhiAck/$entry
      -- 
    convTransposeC_CP_6123_elements(83) <= OrReduce(convTransposeC_CP_6123_elements(75) & convTransposeC_CP_6123_elements(82));
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_2155/merge_stmt_2296_PhiAck/phi_stmt_2297_ack
      -- 
    phi_stmt_2297_ack_7192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2297_ack_0, ack => convTransposeC_CP_6123_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2155/merge_stmt_2296_PhiAck/phi_stmt_2304_ack
      -- 
    phi_stmt_2304_ack_7193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2304_ack_0, ack => convTransposeC_CP_6123_elements(85)); -- 
    -- CP-element group 86:  join  fork  transition  place  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	32 
    -- CP-element group 86: 	33 
    -- CP-element group 86: 	34 
    -- CP-element group 86: 	35 
    -- CP-element group 86:  members (16) 
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2314_update_start_
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2314_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_2155/merge_stmt_2296__exit__
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422__entry__
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2314_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2314_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2314_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2314_Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2319_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2319_update_start_
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2319_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2319_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2319_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/type_cast_2319_Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2155/assign_stmt_2315_to_assign_stmt_2422/$entry
      -- CP-element group 86: 	 branch_block_stmt_2155/merge_stmt_2296_PhiAck/$exit
      -- 
    rr_6730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(86), ack => type_cast_2314_inst_req_0); -- 
    cr_6735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(86), ack => type_cast_2314_inst_req_1); -- 
    rr_6744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(86), ack => type_cast_2319_inst_req_0); -- 
    cr_6749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(86), ack => type_cast_2319_inst_req_1); -- 
    convTransposeC_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6123_elements(84) & convTransposeC_CP_6123_elements(85);
      gj_convTransposeC_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6123_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	59 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Sample/ra
      -- 
    ra_7213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2431_inst_ack_0, ack => convTransposeC_CP_6123_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	59 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Update/ca
      -- 
    ca_7218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2431_inst_ack_1, ack => convTransposeC_CP_6123_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 89: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/$exit
      -- CP-element group 89: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/$exit
      -- CP-element group 89: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_2155/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_req
      -- 
    phi_stmt_2425_req_7219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2425_req_7219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(89), ack => phi_stmt_2425_req_1); -- 
    convTransposeC_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6123_elements(87) & convTransposeC_CP_6123_elements(88);
      gj_convTransposeC_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6123_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  output  delay-element  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	36 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2155/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 90: 	 branch_block_stmt_2155/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2425/$exit
      -- CP-element group 90: 	 branch_block_stmt_2155/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2155/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2429_konst_delay_trans
      -- CP-element group 90: 	 branch_block_stmt_2155/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2425/phi_stmt_2425_req
      -- 
    phi_stmt_2425_req_7230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2425_req_7230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(90), ack => phi_stmt_2425_req_0); -- 
    -- Element group convTransposeC_CP_6123_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => convTransposeC_CP_6123_elements(36), ack => convTransposeC_CP_6123_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  merge  transition  place  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2155/merge_stmt_2424_PhiReqMerge
      -- CP-element group 91: 	 branch_block_stmt_2155/merge_stmt_2424_PhiAck/$entry
      -- 
    convTransposeC_CP_6123_elements(91) <= OrReduce(convTransposeC_CP_6123_elements(90) & convTransposeC_CP_6123_elements(89));
    -- CP-element group 92:  fork  transition  place  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	37 
    -- CP-element group 92: 	38 
    -- CP-element group 92: 	40 
    -- CP-element group 92: 	42 
    -- CP-element group 92: 	44 
    -- CP-element group 92: 	46 
    -- CP-element group 92: 	50 
    -- CP-element group 92: 	52 
    -- CP-element group 92: 	48 
    -- CP-element group 92: 	55 
    -- CP-element group 92: 	56 
    -- CP-element group 92: 	57 
    -- CP-element group 92:  members (45) 
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2478_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2478_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2502_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2441_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530__entry__
      -- CP-element group 92: 	 branch_block_stmt_2155/merge_stmt_2424__exit__
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2471_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2471_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2471_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2478_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2502_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2502_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2441_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2441_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2482_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2441_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2509_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2441_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2441_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2477_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/array_obj_ref_2508_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2509_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/addr_of_2509_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/ptr_deref_2512_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2518_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2518_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2518_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2518_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2518_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2155/assign_stmt_2438_to_assign_stmt_2530/type_cast_2518_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2155/merge_stmt_2424_PhiAck/$exit
      -- CP-element group 92: 	 branch_block_stmt_2155/merge_stmt_2424_PhiAck/phi_stmt_2425_ack
      -- 
    phi_stmt_2425_ack_7235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2425_ack_0, ack => convTransposeC_CP_6123_elements(92)); -- 
    cr_6871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(92), ack => ptr_deref_2482_load_0_req_1); -- 
    req_6826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(92), ack => addr_of_2478_final_reg_req_1); -- 
    cr_6780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(92), ack => type_cast_2471_inst_req_1); -- 
    req_6811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(92), ack => array_obj_ref_2477_index_offset_req_1); -- 
    cr_6890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(92), ack => type_cast_2502_inst_req_1); -- 
    cr_6766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(92), ack => type_cast_2441_inst_req_1); -- 
    rr_6761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(92), ack => type_cast_2441_inst_req_0); -- 
    req_6921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(92), ack => array_obj_ref_2508_index_offset_req_1); -- 
    req_6936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(92), ack => addr_of_2509_final_reg_req_1); -- 
    cr_6986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(92), ack => ptr_deref_2512_store_0_req_1); -- 
    rr_6995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(92), ack => type_cast_2518_inst_req_0); -- 
    cr_7000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6123_elements(92), ack => type_cast_2518_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2384_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2405_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2465_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2496_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_2233_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2233_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom62_2507_resized : std_logic_vector(13 downto 0);
    signal R_idxprom62_2507_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2476_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2476_scaled : std_logic_vector(13 downto 0);
    signal add18_2447 : std_logic_vector(31 downto 0);
    signal add26_2345 : std_logic_vector(31 downto 0);
    signal add37_2360 : std_logic_vector(31 downto 0);
    signal add52_2417 : std_logic_vector(31 downto 0);
    signal add54_2452 : std_logic_vector(31 downto 0);
    signal add67_2525 : std_logic_vector(31 downto 0);
    signal add_2330 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2477_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2477_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2477_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2477_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2477_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2477_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2508_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2508_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2508_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2508_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2508_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2508_root_address : std_logic_vector(13 downto 0);
    signal arrayidx63_2510 : std_logic_vector(31 downto 0);
    signal arrayidx_2479 : std_logic_vector(31 downto 0);
    signal call_2158 : std_logic_vector(15 downto 0);
    signal cmp79_2561 : std_logic_vector(0 downto 0);
    signal cmp87_2587 : std_logic_vector(0 downto 0);
    signal cmp_2530 : std_logic_vector(0 downto 0);
    signal conv10100_2442 : std_logic_vector(31 downto 0);
    signal conv13_2315 : std_logic_vector(31 downto 0);
    signal conv16_2320 : std_logic_vector(31 downto 0);
    signal conv23_2219 : std_logic_vector(31 downto 0);
    signal conv28_2238 : std_logic_vector(31 downto 0);
    signal conv34_2252 : std_logic_vector(31 downto 0);
    signal conv47_2386 : std_logic_vector(31 downto 0);
    signal conv50_2407 : std_logic_vector(31 downto 0);
    signal conv66_2519 : std_logic_vector(31 downto 0);
    signal conv76_2556 : std_logic_vector(31 downto 0);
    signal conv85_2582 : std_logic_vector(31 downto 0);
    signal conv_2181 : std_logic_vector(15 downto 0);
    signal div78_2294 : std_logic_vector(31 downto 0);
    signal div_2177 : std_logic_vector(31 downto 0);
    signal iNsTr_10_2284 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2167 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2189 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2201 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2211 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2227 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2244 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2260 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2272 : std_logic_vector(31 downto 0);
    signal idxprom62_2503 : std_logic_vector(63 downto 0);
    signal idxprom_2472 : std_logic_vector(63 downto 0);
    signal inc83_2565 : std_logic_vector(15 downto 0);
    signal inc83x_xinput_dim0x_x2_2570 : std_logic_vector(15 downto 0);
    signal inc_2551 : std_logic_vector(15 downto 0);
    signal indvar_2425 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2543 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2304 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2297 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2577 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2438 : std_logic_vector(15 downto 0);
    signal mul17_2335 : std_logic_vector(31 downto 0);
    signal mul24_2340 : std_logic_vector(31 downto 0);
    signal mul35_2355 : std_logic_vector(31 downto 0);
    signal mul51_2412 : std_logic_vector(31 downto 0);
    signal mul53_2422 : std_logic_vector(31 downto 0);
    signal mul_2325 : std_logic_vector(31 downto 0);
    signal ptr_deref_2170_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2170_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2170_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2170_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2170_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2192_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2192_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2192_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2192_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2192_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2204_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2204_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2204_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2204_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2204_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2214_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2214_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2214_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2214_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2214_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2230_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2230_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2230_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2230_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2230_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2247_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2247_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2247_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2247_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2247_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2263_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2263_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2263_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2263_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2263_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2275_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2275_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2275_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2275_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2275_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2287_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2287_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2287_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2287_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2287_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2482_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2482_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2482_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2482_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2482_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2512_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2512_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2512_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2512_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2512_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2512_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext101_2398 : std_logic_vector(31 downto 0);
    signal sext103_2458 : std_logic_vector(31 downto 0);
    signal sext104_2489 : std_logic_vector(31 downto 0);
    signal sext_2377 : std_logic_vector(31 downto 0);
    signal shr61_2498 : std_logic_vector(31 downto 0);
    signal shr_2467 : std_logic_vector(31 downto 0);
    signal sub29_2392 : std_logic_vector(31 downto 0);
    signal sub40_2365 : std_logic_vector(31 downto 0);
    signal sub41_2371 : std_logic_vector(31 downto 0);
    signal sub_2350 : std_logic_vector(31 downto 0);
    signal tmp11_2193 : std_logic_vector(31 downto 0);
    signal tmp14_2205 : std_logic_vector(31 downto 0);
    signal tmp22_2215 : std_logic_vector(15 downto 0);
    signal tmp25_2231 : std_logic_vector(31 downto 0);
    signal tmp27_2234 : std_logic_vector(15 downto 0);
    signal tmp33_2248 : std_logic_vector(15 downto 0);
    signal tmp36_2264 : std_logic_vector(31 downto 0);
    signal tmp45_2276 : std_logic_vector(31 downto 0);
    signal tmp48_2288 : std_logic_vector(31 downto 0);
    signal tmp58_2483 : std_logic_vector(63 downto 0);
    signal tmp_2171 : std_logic_vector(31 downto 0);
    signal type_cast_2175_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2292_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2300_wire : std_logic_vector(15 downto 0);
    signal type_cast_2303_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2307_wire : std_logic_vector(15 downto 0);
    signal type_cast_2309_wire : std_logic_vector(15 downto 0);
    signal type_cast_2313_wire : std_logic_vector(31 downto 0);
    signal type_cast_2318_wire : std_logic_vector(31 downto 0);
    signal type_cast_2369_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2375_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2380_wire : std_logic_vector(31 downto 0);
    signal type_cast_2383_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2390_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2396_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2401_wire : std_logic_vector(31 downto 0);
    signal type_cast_2404_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2429_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2431_wire : std_logic_vector(15 downto 0);
    signal type_cast_2436_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2456_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2461_wire : std_logic_vector(31 downto 0);
    signal type_cast_2464_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2470_wire : std_logic_vector(63 downto 0);
    signal type_cast_2487_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2492_wire : std_logic_vector(31 downto 0);
    signal type_cast_2495_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2501_wire : std_logic_vector(63 downto 0);
    signal type_cast_2517_wire : std_logic_vector(31 downto 0);
    signal type_cast_2523_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2541_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2549_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2554_wire : std_logic_vector(31 downto 0);
    signal type_cast_2574_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2580_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_2233_word_address_0 <= "0";
    array_obj_ref_2477_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2477_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2477_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2477_resized_base_address <= "00000000000000";
    array_obj_ref_2508_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2508_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2508_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2508_resized_base_address <= "00000000000000";
    iNsTr_10_2284 <= "00000000000000000000000000000011";
    iNsTr_2_2167 <= "00000000000000000000000000000010";
    iNsTr_3_2189 <= "00000000000000000000000000000100";
    iNsTr_4_2201 <= "00000000000000000000000000000011";
    iNsTr_5_2211 <= "00000000000000000000000000000000";
    iNsTr_6_2227 <= "00000000000000000000000000000011";
    iNsTr_7_2244 <= "00000000000000000000000000000001";
    iNsTr_8_2260 <= "00000000000000000000000000000100";
    iNsTr_9_2272 <= "00000000000000000000000000000100";
    ptr_deref_2170_word_offset_0 <= "0000000";
    ptr_deref_2192_word_offset_0 <= "0000000";
    ptr_deref_2204_word_offset_0 <= "0000000";
    ptr_deref_2214_word_offset_0 <= "0";
    ptr_deref_2230_word_offset_0 <= "0000000";
    ptr_deref_2247_word_offset_0 <= "0";
    ptr_deref_2263_word_offset_0 <= "0000000";
    ptr_deref_2275_word_offset_0 <= "0000000";
    ptr_deref_2287_word_offset_0 <= "0000000";
    ptr_deref_2482_word_offset_0 <= "00000000000000";
    ptr_deref_2512_word_offset_0 <= "00000000000000";
    type_cast_2175_wire_constant <= "00000000000000000000000000000001";
    type_cast_2292_wire_constant <= "00000000000000000000000000000001";
    type_cast_2303_wire_constant <= "0000000000000000";
    type_cast_2369_wire_constant <= "00000000000000000000000000010000";
    type_cast_2375_wire_constant <= "11111111111111110000000000000000";
    type_cast_2383_wire_constant <= "00000000000000000000000000010000";
    type_cast_2390_wire_constant <= "00000000000000000000000000010000";
    type_cast_2396_wire_constant <= "11111111111111110000000000000000";
    type_cast_2404_wire_constant <= "00000000000000000000000000010000";
    type_cast_2429_wire_constant <= "0000000000000000";
    type_cast_2436_wire_constant <= "0000000000000100";
    type_cast_2456_wire_constant <= "00000000000000000000000000010000";
    type_cast_2464_wire_constant <= "00000000000000000000000000010010";
    type_cast_2487_wire_constant <= "00000000000000000000000000010000";
    type_cast_2495_wire_constant <= "00000000000000000000000000010010";
    type_cast_2523_wire_constant <= "00000000000000000000000000000100";
    type_cast_2541_wire_constant <= "0000000000000001";
    type_cast_2549_wire_constant <= "0000000000000001";
    type_cast_2574_wire_constant <= "0000000000000000";
    phi_stmt_2297: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2300_wire & type_cast_2303_wire_constant;
      req <= phi_stmt_2297_req_0 & phi_stmt_2297_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2297",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2297_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2297,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2297
    phi_stmt_2304: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2307_wire & type_cast_2309_wire;
      req <= phi_stmt_2304_req_0 & phi_stmt_2304_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2304",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2304_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2304,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2304
    phi_stmt_2425: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2429_wire_constant & type_cast_2431_wire;
      req <= phi_stmt_2425_req_0 & phi_stmt_2425_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2425",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2425_ack_0,
          idata => idata,
          odata => indvar_2425,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2425
    -- flow-through select operator MUX_2576_inst
    input_dim1x_x2_2577 <= type_cast_2574_wire_constant when (cmp79_2561(0) /=  '0') else inc_2551;
    addr_of_2478_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2478_final_reg_req_0;
      addr_of_2478_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2478_final_reg_req_1;
      addr_of_2478_final_reg_ack_1<= rack(0);
      addr_of_2478_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2478_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2477_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2479,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2509_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2509_final_reg_req_0;
      addr_of_2509_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2509_final_reg_req_1;
      addr_of_2509_final_reg_ack_1<= rack(0);
      addr_of_2509_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2509_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2508_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx63_2510,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2180_inst_req_0;
      type_cast_2180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2180_inst_req_1;
      type_cast_2180_inst_ack_1<= rack(0);
      type_cast_2180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2180_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2177,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2181,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2218_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2218_inst_req_0;
      type_cast_2218_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2218_inst_req_1;
      type_cast_2218_inst_ack_1<= rack(0);
      type_cast_2218_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2218_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp22_2215,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_2219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2237_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2237_inst_req_0;
      type_cast_2237_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2237_inst_req_1;
      type_cast_2237_inst_ack_1<= rack(0);
      type_cast_2237_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2237_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp27_2234,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv28_2238,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2251_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2251_inst_req_0;
      type_cast_2251_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2251_inst_req_1;
      type_cast_2251_inst_ack_1<= rack(0);
      type_cast_2251_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2251_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp33_2248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv34_2252,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2300_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2300_inst_req_0;
      type_cast_2300_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2300_inst_req_1;
      type_cast_2300_inst_ack_1<= rack(0);
      type_cast_2300_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2300_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2577,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2300_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2307_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2307_inst_req_0;
      type_cast_2307_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2307_inst_req_1;
      type_cast_2307_inst_ack_1<= rack(0);
      type_cast_2307_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2307_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc83x_xinput_dim0x_x2_2570,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2307_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2309_inst_req_0;
      type_cast_2309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2309_inst_req_1;
      type_cast_2309_inst_ack_1<= rack(0);
      type_cast_2309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_2181,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2309_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2314_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2314_inst_req_0;
      type_cast_2314_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2314_inst_req_1;
      type_cast_2314_inst_ack_1<= rack(0);
      type_cast_2314_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2314_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2313_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13_2315,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2319_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2319_inst_req_0;
      type_cast_2319_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2319_inst_req_1;
      type_cast_2319_inst_ack_1<= rack(0);
      type_cast_2319_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2319_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2318_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_2320,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2380_inst
    process(sext_2377) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2377(31 downto 0);
      type_cast_2380_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2385_inst
    process(ASHR_i32_i32_2384_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2384_wire(31 downto 0);
      conv47_2386 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2401_inst
    process(sext101_2398) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext101_2398(31 downto 0);
      type_cast_2401_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2406_inst
    process(ASHR_i32_i32_2405_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2405_wire(31 downto 0);
      conv50_2407 <= tmp_var; -- 
    end process;
    type_cast_2431_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2431_inst_req_0;
      type_cast_2431_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2431_inst_req_1;
      type_cast_2431_inst_ack_1<= rack(0);
      type_cast_2431_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2431_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2543,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2431_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2441_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2441_inst_req_0;
      type_cast_2441_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2441_inst_req_1;
      type_cast_2441_inst_ack_1<= rack(0);
      type_cast_2441_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2441_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2438,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10100_2442,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2461_inst
    process(sext103_2458) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext103_2458(31 downto 0);
      type_cast_2461_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2466_inst
    process(ASHR_i32_i32_2465_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2465_wire(31 downto 0);
      shr_2467 <= tmp_var; -- 
    end process;
    type_cast_2471_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2471_inst_req_0;
      type_cast_2471_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2471_inst_req_1;
      type_cast_2471_inst_ack_1<= rack(0);
      type_cast_2471_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2471_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2470_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2472,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2492_inst
    process(sext104_2489) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext104_2489(31 downto 0);
      type_cast_2492_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2497_inst
    process(ASHR_i32_i32_2496_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2496_wire(31 downto 0);
      shr61_2498 <= tmp_var; -- 
    end process;
    type_cast_2502_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2502_inst_req_0;
      type_cast_2502_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2502_inst_req_1;
      type_cast_2502_inst_ack_1<= rack(0);
      type_cast_2502_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2502_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2501_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom62_2503,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2518_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2518_inst_req_0;
      type_cast_2518_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2518_inst_req_1;
      type_cast_2518_inst_ack_1<= rack(0);
      type_cast_2518_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2518_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2517_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_2519,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2555_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2555_inst_req_0;
      type_cast_2555_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2555_inst_req_1;
      type_cast_2555_inst_ack_1<= rack(0);
      type_cast_2555_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2555_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2554_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_2556,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2564_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2564_inst_req_0;
      type_cast_2564_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2564_inst_req_1;
      type_cast_2564_inst_ack_1<= rack(0);
      type_cast_2564_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2564_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp79_2561,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc83_2565,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2581_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2581_inst_req_0;
      type_cast_2581_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2581_inst_req_1;
      type_cast_2581_inst_ack_1<= rack(0);
      type_cast_2581_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2581_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2580_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_2582,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2233_gather_scatter
    process(LOAD_padding_2233_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2233_data_0;
      ov(15 downto 0) := iv;
      tmp27_2234 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2477_index_1_rename
    process(R_idxprom_2476_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2476_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2476_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2477_index_1_resize
    process(idxprom_2472) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2472;
      ov := iv(13 downto 0);
      R_idxprom_2476_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2477_root_address_inst
    process(array_obj_ref_2477_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2477_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2477_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2508_index_1_rename
    process(R_idxprom62_2507_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom62_2507_resized;
      ov(13 downto 0) := iv;
      R_idxprom62_2507_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2508_index_1_resize
    process(idxprom62_2503) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom62_2503;
      ov := iv(13 downto 0);
      R_idxprom62_2507_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2508_root_address_inst
    process(array_obj_ref_2508_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2508_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2508_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2170_addr_0
    process(ptr_deref_2170_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2170_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2170_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2170_base_resize
    process(iNsTr_2_2167) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2167;
      ov := iv(6 downto 0);
      ptr_deref_2170_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2170_gather_scatter
    process(ptr_deref_2170_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2170_data_0;
      ov(31 downto 0) := iv;
      tmp_2171 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2170_root_address_inst
    process(ptr_deref_2170_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2170_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2170_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2192_addr_0
    process(ptr_deref_2192_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2192_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2192_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2192_base_resize
    process(iNsTr_3_2189) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2189;
      ov := iv(6 downto 0);
      ptr_deref_2192_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2192_gather_scatter
    process(ptr_deref_2192_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2192_data_0;
      ov(31 downto 0) := iv;
      tmp11_2193 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2192_root_address_inst
    process(ptr_deref_2192_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2192_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2192_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2204_addr_0
    process(ptr_deref_2204_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2204_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2204_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2204_base_resize
    process(iNsTr_4_2201) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2201;
      ov := iv(6 downto 0);
      ptr_deref_2204_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2204_gather_scatter
    process(ptr_deref_2204_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2204_data_0;
      ov(31 downto 0) := iv;
      tmp14_2205 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2204_root_address_inst
    process(ptr_deref_2204_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2204_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2204_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2214_addr_0
    process(ptr_deref_2214_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2214_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2214_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2214_base_resize
    process(iNsTr_5_2211) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2211;
      ov := iv(0 downto 0);
      ptr_deref_2214_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2214_gather_scatter
    process(ptr_deref_2214_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2214_data_0;
      ov(15 downto 0) := iv;
      tmp22_2215 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2214_root_address_inst
    process(ptr_deref_2214_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2214_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2214_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2230_addr_0
    process(ptr_deref_2230_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2230_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2230_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2230_base_resize
    process(iNsTr_6_2227) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2227;
      ov := iv(6 downto 0);
      ptr_deref_2230_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2230_gather_scatter
    process(ptr_deref_2230_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2230_data_0;
      ov(31 downto 0) := iv;
      tmp25_2231 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2230_root_address_inst
    process(ptr_deref_2230_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2230_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2230_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2247_addr_0
    process(ptr_deref_2247_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2247_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2247_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2247_base_resize
    process(iNsTr_7_2244) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2244;
      ov := iv(0 downto 0);
      ptr_deref_2247_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2247_gather_scatter
    process(ptr_deref_2247_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2247_data_0;
      ov(15 downto 0) := iv;
      tmp33_2248 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2247_root_address_inst
    process(ptr_deref_2247_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2247_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2247_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2263_addr_0
    process(ptr_deref_2263_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2263_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2263_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2263_base_resize
    process(iNsTr_8_2260) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2260;
      ov := iv(6 downto 0);
      ptr_deref_2263_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2263_gather_scatter
    process(ptr_deref_2263_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2263_data_0;
      ov(31 downto 0) := iv;
      tmp36_2264 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2263_root_address_inst
    process(ptr_deref_2263_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2263_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2263_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2275_addr_0
    process(ptr_deref_2275_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2275_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2275_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2275_base_resize
    process(iNsTr_9_2272) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2272;
      ov := iv(6 downto 0);
      ptr_deref_2275_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2275_gather_scatter
    process(ptr_deref_2275_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2275_data_0;
      ov(31 downto 0) := iv;
      tmp45_2276 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2275_root_address_inst
    process(ptr_deref_2275_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2275_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2275_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2287_addr_0
    process(ptr_deref_2287_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2287_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2287_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2287_base_resize
    process(iNsTr_10_2284) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2284;
      ov := iv(6 downto 0);
      ptr_deref_2287_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2287_gather_scatter
    process(ptr_deref_2287_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2287_data_0;
      ov(31 downto 0) := iv;
      tmp48_2288 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2287_root_address_inst
    process(ptr_deref_2287_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2287_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2287_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2482_addr_0
    process(ptr_deref_2482_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2482_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2482_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2482_base_resize
    process(arrayidx_2479) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2479;
      ov := iv(13 downto 0);
      ptr_deref_2482_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2482_gather_scatter
    process(ptr_deref_2482_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2482_data_0;
      ov(63 downto 0) := iv;
      tmp58_2483 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2482_root_address_inst
    process(ptr_deref_2482_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2482_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2482_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2512_addr_0
    process(ptr_deref_2512_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2512_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2512_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2512_base_resize
    process(arrayidx63_2510) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx63_2510;
      ov := iv(13 downto 0);
      ptr_deref_2512_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2512_gather_scatter
    process(tmp58_2483) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp58_2483;
      ov(63 downto 0) := iv;
      ptr_deref_2512_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2512_root_address_inst
    process(ptr_deref_2512_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2512_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2512_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2531_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2530;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2531_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2531_branch_req_0,
          ack0 => if_stmt_2531_branch_ack_0,
          ack1 => if_stmt_2531_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2588_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp87_2587;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2588_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2588_branch_req_0,
          ack0 => if_stmt_2588_branch_ack_0,
          ack1 => if_stmt_2588_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2542_inst
    process(indvar_2425) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2425, type_cast_2541_wire_constant, tmp_var);
      indvarx_xnext_2543 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2550_inst
    process(input_dim1x_x1x_xph_2297) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2297, type_cast_2549_wire_constant, tmp_var);
      inc_2551 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2569_inst
    process(inc83_2565, input_dim0x_x2x_xph_2304) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc83_2565, input_dim0x_x2x_xph_2304, tmp_var);
      inc83x_xinput_dim0x_x2_2570 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2329_inst
    process(mul_2325, conv13_2315) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_2325, conv13_2315, tmp_var);
      add_2330 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2344_inst
    process(mul24_2340, tmp25_2231) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul24_2340, tmp25_2231, tmp_var);
      add26_2345 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2359_inst
    process(mul35_2355, tmp36_2264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul35_2355, tmp36_2264, tmp_var);
      add37_2360 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2376_inst
    process(sub41_2371) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub41_2371, type_cast_2375_wire_constant, tmp_var);
      sext_2377 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2397_inst
    process(sub29_2392) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub29_2392, type_cast_2396_wire_constant, tmp_var);
      sext101_2398 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2416_inst
    process(conv47_2386, mul51_2412) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv47_2386, mul51_2412, tmp_var);
      add52_2417 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2446_inst
    process(mul17_2335, conv10100_2442) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul17_2335, conv10100_2442, tmp_var);
      add18_2447 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2451_inst
    process(mul53_2422, conv10100_2442) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul53_2422, conv10100_2442, tmp_var);
      add54_2452 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2524_inst
    process(conv66_2519) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv66_2519, type_cast_2523_wire_constant, tmp_var);
      add67_2525 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2384_inst
    process(type_cast_2380_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2380_wire, type_cast_2383_wire_constant, tmp_var);
      ASHR_i32_i32_2384_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2405_inst
    process(type_cast_2401_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2401_wire, type_cast_2404_wire_constant, tmp_var);
      ASHR_i32_i32_2405_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2465_inst
    process(type_cast_2461_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2461_wire, type_cast_2464_wire_constant, tmp_var);
      ASHR_i32_i32_2465_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2496_inst
    process(type_cast_2492_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2492_wire, type_cast_2495_wire_constant, tmp_var);
      ASHR_i32_i32_2496_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2560_inst
    process(conv76_2556, div78_2294) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv76_2556, div78_2294, tmp_var);
      cmp79_2561 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2586_inst
    process(conv85_2582, tmp_2171) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv85_2582, tmp_2171, tmp_var);
      cmp87_2587 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2176_inst
    process(tmp_2171) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2171, type_cast_2175_wire_constant, tmp_var);
      div_2177 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2293_inst
    process(tmp14_2205) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_2205, type_cast_2292_wire_constant, tmp_var);
      div78_2294 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2437_inst
    process(indvar_2425) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2425, type_cast_2436_wire_constant, tmp_var);
      input_dim2x_x1_2438 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2324_inst
    process(tmp14_2205, conv16_2320) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_2205, conv16_2320, tmp_var);
      mul_2325 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2334_inst
    process(add_2330, tmp11_2193) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_2330, tmp11_2193, tmp_var);
      mul17_2335 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2339_inst
    process(conv23_2219, conv16_2320) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv23_2219, conv16_2320, tmp_var);
      mul24_2340 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2354_inst
    process(conv34_2252, conv13_2315) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv34_2252, conv13_2315, tmp_var);
      mul35_2355 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2411_inst
    process(tmp48_2288, conv50_2407) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp48_2288, conv50_2407, tmp_var);
      mul51_2412 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2421_inst
    process(add52_2417, tmp45_2276) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add52_2417, tmp45_2276, tmp_var);
      mul53_2422 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2370_inst
    process(sub40_2365) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub40_2365, type_cast_2369_wire_constant, tmp_var);
      sub41_2371 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2391_inst
    process(sub_2350) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2350, type_cast_2390_wire_constant, tmp_var);
      sub29_2392 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2457_inst
    process(add18_2447) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add18_2447, type_cast_2456_wire_constant, tmp_var);
      sext103_2458 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2488_inst
    process(add54_2452) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add54_2452, type_cast_2487_wire_constant, tmp_var);
      sext104_2489 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2349_inst
    process(add26_2345, conv28_2238) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add26_2345, conv28_2238, tmp_var);
      sub_2350 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2364_inst
    process(add37_2360, conv28_2238) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add37_2360, conv28_2238, tmp_var);
      sub40_2365 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2529_inst
    process(add67_2525, tmp11_2193) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add67_2525, tmp11_2193, tmp_var);
      cmp_2530 <= tmp_var; --
    end process;
    -- shared split operator group (34) : array_obj_ref_2477_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2476_scaled;
      array_obj_ref_2477_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2477_index_offset_req_0;
      array_obj_ref_2477_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2477_index_offset_req_1;
      array_obj_ref_2477_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_2508_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom62_2507_scaled;
      array_obj_ref_2508_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2508_index_offset_req_0;
      array_obj_ref_2508_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2508_index_offset_req_1;
      array_obj_ref_2508_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- unary operator type_cast_2313_inst
    process(input_dim1x_x1x_xph_2297) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_2297, tmp_var);
      type_cast_2313_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2318_inst
    process(input_dim0x_x2x_xph_2304) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_2304, tmp_var);
      type_cast_2318_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2470_inst
    process(shr_2467) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2467, tmp_var);
      type_cast_2470_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2501_inst
    process(shr61_2498) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr61_2498, tmp_var);
      type_cast_2501_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2517_inst
    process(input_dim2x_x1_2438) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2438, tmp_var);
      type_cast_2517_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2554_inst
    process(inc_2551) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2551, tmp_var);
      type_cast_2554_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2580_inst
    process(inc83x_xinput_dim0x_x2_2570) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc83x_xinput_dim0x_x2_2570, tmp_var);
      type_cast_2580_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_2233_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2233_load_0_req_0;
      LOAD_padding_2233_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2233_load_0_req_1;
      LOAD_padding_2233_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2233_word_address_0;
      LOAD_padding_2233_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2204_load_0 ptr_deref_2192_load_0 ptr_deref_2170_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2204_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2192_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2170_load_0_req_0;
      ptr_deref_2204_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2192_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2170_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2204_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2192_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2170_load_0_req_1;
      ptr_deref_2204_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2192_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2170_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2204_word_address_0 & ptr_deref_2192_word_address_0 & ptr_deref_2170_word_address_0;
      ptr_deref_2204_data_0 <= data_out(95 downto 64);
      ptr_deref_2192_data_0 <= data_out(63 downto 32);
      ptr_deref_2170_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2247_load_0 ptr_deref_2214_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2247_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2214_load_0_req_0;
      ptr_deref_2247_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2214_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2247_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2214_load_0_req_1;
      ptr_deref_2247_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2214_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2247_word_address_0 & ptr_deref_2214_word_address_0;
      ptr_deref_2247_data_0 <= data_out(31 downto 16);
      ptr_deref_2214_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2263_load_0 ptr_deref_2230_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2263_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2230_load_0_req_0;
      ptr_deref_2263_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2230_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2263_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2230_load_0_req_1;
      ptr_deref_2263_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2230_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2263_word_address_0 & ptr_deref_2230_word_address_0;
      ptr_deref_2263_data_0 <= data_out(63 downto 32);
      ptr_deref_2230_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2275_load_0 ptr_deref_2287_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2275_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2287_load_0_req_0;
      ptr_deref_2275_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2287_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2275_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2287_load_0_req_1;
      ptr_deref_2275_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2287_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2275_word_address_0 & ptr_deref_2287_word_address_0;
      ptr_deref_2275_data_0 <= data_out(63 downto 32);
      ptr_deref_2287_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2482_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2482_load_0_req_0;
      ptr_deref_2482_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2482_load_0_req_1;
      ptr_deref_2482_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2482_word_address_0;
      ptr_deref_2482_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2512_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2512_store_0_req_0;
      ptr_deref_2512_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2512_store_0_req_1;
      ptr_deref_2512_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2512_word_address_0;
      data_in <= ptr_deref_2512_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2157_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_start_2157_inst_req_0;
      RPIPE_Block2_start_2157_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_start_2157_inst_req_1;
      RPIPE_Block2_start_2157_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2158 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2596_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2596_inst_req_0;
      WPIPE_Block2_done_2596_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2596_inst_req_1;
      WPIPE_Block2_done_2596_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2158;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_7276_start: Boolean;
  signal convTransposeD_CP_7276_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_2619_load_0_ack_0 : boolean;
  signal ptr_deref_2641_load_0_ack_0 : boolean;
  signal ptr_deref_2641_load_0_ack_1 : boolean;
  signal ptr_deref_2641_load_0_req_1 : boolean;
  signal ptr_deref_2641_load_0_req_0 : boolean;
  signal ptr_deref_2619_load_0_ack_1 : boolean;
  signal type_cast_2651_inst_ack_0 : boolean;
  signal type_cast_2677_inst_req_1 : boolean;
  signal type_cast_2629_inst_req_1 : boolean;
  signal type_cast_2629_inst_ack_1 : boolean;
  signal type_cast_2651_inst_req_0 : boolean;
  signal type_cast_3048_inst_ack_1 : boolean;
  signal ptr_deref_2689_load_0_req_1 : boolean;
  signal ptr_deref_2689_load_0_ack_1 : boolean;
  signal type_cast_3048_inst_req_1 : boolean;
  signal type_cast_2651_inst_ack_1 : boolean;
  signal LOAD_padding_2692_load_0_req_0 : boolean;
  signal LOAD_padding_2692_load_0_ack_0 : boolean;
  signal type_cast_2629_inst_ack_0 : boolean;
  signal type_cast_2629_inst_req_0 : boolean;
  signal ptr_deref_2689_load_0_req_0 : boolean;
  signal ptr_deref_2673_load_0_req_1 : boolean;
  signal ptr_deref_2673_load_0_ack_1 : boolean;
  signal ptr_deref_2663_load_0_req_0 : boolean;
  signal ptr_deref_2663_load_0_ack_0 : boolean;
  signal type_cast_2677_inst_ack_1 : boolean;
  signal ptr_deref_2673_load_0_req_0 : boolean;
  signal ptr_deref_2619_load_0_req_0 : boolean;
  signal ptr_deref_2663_load_0_req_1 : boolean;
  signal ptr_deref_2663_load_0_ack_1 : boolean;
  signal ptr_deref_2673_load_0_ack_0 : boolean;
  signal ptr_deref_2689_load_0_ack_0 : boolean;
  signal ptr_deref_2619_load_0_req_1 : boolean;
  signal type_cast_2677_inst_req_0 : boolean;
  signal type_cast_2677_inst_ack_0 : boolean;
  signal type_cast_2696_inst_ack_0 : boolean;
  signal type_cast_2696_inst_req_1 : boolean;
  signal type_cast_2696_inst_ack_1 : boolean;
  signal type_cast_3048_inst_ack_0 : boolean;
  signal LOAD_padding_2692_load_0_req_1 : boolean;
  signal LOAD_padding_2692_load_0_ack_1 : boolean;
  signal phi_stmt_3039_req_0 : boolean;
  signal type_cast_2696_inst_req_0 : boolean;
  signal type_cast_2651_inst_req_1 : boolean;
  signal phi_stmt_3045_req_0 : boolean;
  signal type_cast_3042_inst_req_0 : boolean;
  signal type_cast_3042_inst_ack_0 : boolean;
  signal type_cast_3042_inst_req_1 : boolean;
  signal type_cast_3042_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2606_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2606_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2606_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2606_inst_ack_1 : boolean;
  signal ptr_deref_2706_load_0_req_0 : boolean;
  signal ptr_deref_2706_load_0_ack_0 : boolean;
  signal ptr_deref_2706_load_0_req_1 : boolean;
  signal ptr_deref_2706_load_0_ack_1 : boolean;
  signal type_cast_2710_inst_req_0 : boolean;
  signal type_cast_2710_inst_ack_0 : boolean;
  signal type_cast_2710_inst_req_1 : boolean;
  signal type_cast_2710_inst_ack_1 : boolean;
  signal ptr_deref_2722_load_0_req_0 : boolean;
  signal ptr_deref_2722_load_0_ack_0 : boolean;
  signal ptr_deref_2722_load_0_req_1 : boolean;
  signal ptr_deref_2722_load_0_ack_1 : boolean;
  signal ptr_deref_2734_load_0_req_0 : boolean;
  signal ptr_deref_2734_load_0_ack_0 : boolean;
  signal ptr_deref_2734_load_0_req_1 : boolean;
  signal ptr_deref_2734_load_0_ack_1 : boolean;
  signal ptr_deref_2746_load_0_req_0 : boolean;
  signal ptr_deref_2746_load_0_ack_0 : boolean;
  signal ptr_deref_2746_load_0_req_1 : boolean;
  signal ptr_deref_2746_load_0_ack_1 : boolean;
  signal type_cast_2766_inst_req_0 : boolean;
  signal type_cast_2766_inst_ack_0 : boolean;
  signal type_cast_2766_inst_req_1 : boolean;
  signal type_cast_2766_inst_ack_1 : boolean;
  signal type_cast_2771_inst_req_0 : boolean;
  signal type_cast_2771_inst_ack_0 : boolean;
  signal type_cast_2771_inst_req_1 : boolean;
  signal type_cast_2771_inst_ack_1 : boolean;
  signal type_cast_2893_inst_req_0 : boolean;
  signal type_cast_2893_inst_ack_0 : boolean;
  signal type_cast_2893_inst_req_1 : boolean;
  signal type_cast_2893_inst_ack_1 : boolean;
  signal type_cast_2923_inst_req_0 : boolean;
  signal type_cast_2923_inst_ack_0 : boolean;
  signal type_cast_3048_inst_req_0 : boolean;
  signal type_cast_2923_inst_req_1 : boolean;
  signal type_cast_2923_inst_ack_1 : boolean;
  signal array_obj_ref_2929_index_offset_req_0 : boolean;
  signal array_obj_ref_2929_index_offset_ack_0 : boolean;
  signal array_obj_ref_2929_index_offset_req_1 : boolean;
  signal array_obj_ref_2929_index_offset_ack_1 : boolean;
  signal phi_stmt_3045_ack_0 : boolean;
  signal addr_of_2930_final_reg_req_0 : boolean;
  signal addr_of_2930_final_reg_ack_0 : boolean;
  signal addr_of_2930_final_reg_req_1 : boolean;
  signal addr_of_2930_final_reg_ack_1 : boolean;
  signal ptr_deref_2934_load_0_req_0 : boolean;
  signal ptr_deref_2934_load_0_ack_0 : boolean;
  signal ptr_deref_2934_load_0_req_1 : boolean;
  signal ptr_deref_2934_load_0_ack_1 : boolean;
  signal type_cast_2954_inst_req_0 : boolean;
  signal type_cast_2954_inst_ack_0 : boolean;
  signal type_cast_2954_inst_req_1 : boolean;
  signal type_cast_2954_inst_ack_1 : boolean;
  signal array_obj_ref_2960_index_offset_req_0 : boolean;
  signal array_obj_ref_2960_index_offset_ack_0 : boolean;
  signal phi_stmt_3039_ack_0 : boolean;
  signal array_obj_ref_2960_index_offset_req_1 : boolean;
  signal array_obj_ref_2960_index_offset_ack_1 : boolean;
  signal addr_of_2961_final_reg_req_0 : boolean;
  signal addr_of_2961_final_reg_ack_0 : boolean;
  signal addr_of_2961_final_reg_req_1 : boolean;
  signal addr_of_2961_final_reg_ack_1 : boolean;
  signal ptr_deref_2964_store_0_req_0 : boolean;
  signal ptr_deref_2964_store_0_ack_0 : boolean;
  signal ptr_deref_2964_store_0_req_1 : boolean;
  signal ptr_deref_2964_store_0_ack_1 : boolean;
  signal type_cast_2970_inst_req_0 : boolean;
  signal type_cast_2970_inst_ack_0 : boolean;
  signal type_cast_2970_inst_req_1 : boolean;
  signal type_cast_2970_inst_ack_1 : boolean;
  signal if_stmt_2983_branch_req_0 : boolean;
  signal if_stmt_2983_branch_ack_1 : boolean;
  signal if_stmt_2983_branch_ack_0 : boolean;
  signal type_cast_3007_inst_req_0 : boolean;
  signal type_cast_3007_inst_ack_0 : boolean;
  signal type_cast_3007_inst_req_1 : boolean;
  signal type_cast_3007_inst_ack_1 : boolean;
  signal if_stmt_3014_branch_req_0 : boolean;
  signal if_stmt_3014_branch_ack_1 : boolean;
  signal if_stmt_3014_branch_ack_0 : boolean;
  signal type_cast_3035_inst_req_0 : boolean;
  signal type_cast_3035_inst_ack_0 : boolean;
  signal type_cast_3035_inst_req_1 : boolean;
  signal type_cast_3035_inst_ack_1 : boolean;
  signal type_cast_3055_inst_req_0 : boolean;
  signal type_cast_3055_inst_ack_0 : boolean;
  signal type_cast_3055_inst_req_1 : boolean;
  signal type_cast_3055_inst_ack_1 : boolean;
  signal if_stmt_3062_branch_req_0 : boolean;
  signal if_stmt_3062_branch_ack_1 : boolean;
  signal if_stmt_3062_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_3070_inst_req_0 : boolean;
  signal WPIPE_Block3_done_3070_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_3070_inst_req_1 : boolean;
  signal WPIPE_Block3_done_3070_inst_ack_1 : boolean;
  signal type_cast_2753_inst_req_0 : boolean;
  signal type_cast_2753_inst_ack_0 : boolean;
  signal type_cast_2753_inst_req_1 : boolean;
  signal type_cast_2753_inst_ack_1 : boolean;
  signal phi_stmt_2750_req_0 : boolean;
  signal type_cast_2759_inst_req_0 : boolean;
  signal type_cast_2759_inst_ack_0 : boolean;
  signal type_cast_2759_inst_req_1 : boolean;
  signal type_cast_2759_inst_ack_1 : boolean;
  signal phi_stmt_2756_req_0 : boolean;
  signal type_cast_2755_inst_req_0 : boolean;
  signal type_cast_2755_inst_ack_0 : boolean;
  signal type_cast_2755_inst_req_1 : boolean;
  signal type_cast_2755_inst_ack_1 : boolean;
  signal phi_stmt_2750_req_1 : boolean;
  signal type_cast_2761_inst_req_0 : boolean;
  signal type_cast_2761_inst_ack_0 : boolean;
  signal type_cast_2761_inst_req_1 : boolean;
  signal type_cast_2761_inst_ack_1 : boolean;
  signal phi_stmt_2756_req_1 : boolean;
  signal phi_stmt_2750_ack_0 : boolean;
  signal phi_stmt_2756_ack_0 : boolean;
  signal type_cast_2883_inst_req_0 : boolean;
  signal type_cast_2883_inst_ack_0 : boolean;
  signal type_cast_2883_inst_req_1 : boolean;
  signal type_cast_2883_inst_ack_1 : boolean;
  signal phi_stmt_2877_req_1 : boolean;
  signal phi_stmt_2877_req_0 : boolean;
  signal phi_stmt_2877_ack_0 : boolean;
  signal type_cast_3044_inst_req_0 : boolean;
  signal type_cast_3044_inst_ack_0 : boolean;
  signal type_cast_3044_inst_req_1 : boolean;
  signal type_cast_3044_inst_ack_1 : boolean;
  signal phi_stmt_3039_req_1 : boolean;
  signal type_cast_3050_inst_req_0 : boolean;
  signal type_cast_3050_inst_ack_0 : boolean;
  signal type_cast_3050_inst_req_1 : boolean;
  signal type_cast_3050_inst_ack_1 : boolean;
  signal phi_stmt_3045_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_7276_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_7276_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_7276_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_7276_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_7276: Block -- control-path 
    signal convTransposeD_CP_7276_elements: BooleanArray(116 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_7276_elements(0) <= convTransposeD_CP_7276_start;
    convTransposeD_CP_7276_symbol <= convTransposeD_CP_7276_elements(74);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2604/$entry
      -- CP-element group 0: 	 branch_block_stmt_2604/branch_block_stmt_2604__entry__
      -- CP-element group 0: 	 branch_block_stmt_2604/assign_stmt_2607__entry__
      -- CP-element group 0: 	 branch_block_stmt_2604/assign_stmt_2607/$entry
      -- CP-element group 0: 	 branch_block_stmt_2604/assign_stmt_2607/RPIPE_Block3_start_2606_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2604/assign_stmt_2607/RPIPE_Block3_start_2606_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2604/assign_stmt_2607/RPIPE_Block3_start_2606_Sample/rr
      -- 
    rr_7334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(0), ack => RPIPE_Block3_start_2606_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2604/assign_stmt_2607/RPIPE_Block3_start_2606_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2604/assign_stmt_2607/RPIPE_Block3_start_2606_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2604/assign_stmt_2607/RPIPE_Block3_start_2606_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2604/assign_stmt_2607/RPIPE_Block3_start_2606_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2604/assign_stmt_2607/RPIPE_Block3_start_2606_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2604/assign_stmt_2607/RPIPE_Block3_start_2606_Update/cr
      -- 
    ra_7335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2606_inst_ack_0, ack => convTransposeD_CP_7276_elements(1)); -- 
    cr_7339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(1), ack => RPIPE_Block3_start_2606_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	32 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	31 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2:  members (268) 
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2651_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2677_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2677_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2629_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2629_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2651_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2677_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2696_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2696_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2696_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2629_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2651_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2607__exit__
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747__entry__
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2607/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2607/RPIPE_Block3_start_2606_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2607/RPIPE_Block3_start_2606_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2607/RPIPE_Block3_start_2606_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2710_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2710_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2710_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Update/word_access_complete/word_0/cr
      -- 
    ca_7340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2606_inst_ack_1, ack => convTransposeD_CP_7276_elements(2)); -- 
    cr_7451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2641_load_0_req_1); -- 
    rr_7440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2641_load_0_req_0); -- 
    cr_7584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => type_cast_2677_inst_req_1); -- 
    cr_7406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => type_cast_2629_inst_req_1); -- 
    cr_7629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2689_load_0_req_1); -- 
    rr_7651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => LOAD_padding_2692_load_0_req_0); -- 
    rr_7618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2689_load_0_req_0); -- 
    cr_7565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2673_load_0_req_1); -- 
    rr_7504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2663_load_0_req_0); -- 
    rr_7554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2673_load_0_req_0); -- 
    rr_7376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2619_load_0_req_0); -- 
    cr_7515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2663_load_0_req_1); -- 
    cr_7387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2619_load_0_req_1); -- 
    cr_7681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => type_cast_2696_inst_req_1); -- 
    cr_7662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => LOAD_padding_2692_load_0_req_1); -- 
    cr_7470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => type_cast_2651_inst_req_1); -- 
    rr_7715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2706_load_0_req_0); -- 
    cr_7726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2706_load_0_req_1); -- 
    cr_7745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => type_cast_2710_inst_req_1); -- 
    rr_7779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2722_load_0_req_0); -- 
    cr_7790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2722_load_0_req_1); -- 
    rr_7829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2734_load_0_req_0); -- 
    cr_7840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2734_load_0_req_1); -- 
    rr_7879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2746_load_0_req_0); -- 
    cr_7890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(2), ack => ptr_deref_2746_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_sample_completed_
      -- 
    ra_7377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2619_load_0_ack_0, ack => convTransposeD_CP_7276_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Update/ptr_deref_2619_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Update/ptr_deref_2619_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Update/ptr_deref_2619_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2629_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_Update/ptr_deref_2619_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2629_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2629_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2619_update_completed_
      -- 
    ca_7388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2619_load_0_ack_1, ack => convTransposeD_CP_7276_elements(4)); -- 
    rr_7401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(4), ack => type_cast_2629_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2629_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2629_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2629_sample_completed_
      -- 
    ra_7402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2629_inst_ack_0, ack => convTransposeD_CP_7276_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	33 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2629_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2629_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2629_update_completed_
      -- 
    ca_7407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2629_inst_ack_1, ack => convTransposeD_CP_7276_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Sample/word_access_start/$exit
      -- 
    ra_7441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2641_load_0_ack_0, ack => convTransposeD_CP_7276_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Update/ptr_deref_2641_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Update/ptr_deref_2641_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Update/ptr_deref_2641_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2651_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2651_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2641_Update/ptr_deref_2641_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2651_Sample/$entry
      -- 
    ca_7452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2641_load_0_ack_1, ack => convTransposeD_CP_7276_elements(8)); -- 
    rr_7465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(8), ack => type_cast_2651_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2651_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2651_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2651_Sample/$exit
      -- 
    ra_7466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2651_inst_ack_0, ack => convTransposeD_CP_7276_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	33 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2651_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2651_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2651_Update/ca
      -- 
    ca_7471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2651_inst_ack_1, ack => convTransposeD_CP_7276_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Sample/word_access_start/word_0/ra
      -- CP-element group 11: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_sample_completed_
      -- 
    ra_7505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2663_load_0_ack_0, ack => convTransposeD_CP_7276_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	33 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Update/ptr_deref_2663_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Update/ptr_deref_2663_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Update/ptr_deref_2663_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Update/ptr_deref_2663_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2663_Update/$exit
      -- 
    ca_7516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2663_load_0_ack_1, ack => convTransposeD_CP_7276_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Sample/word_access_start/word_0/ra
      -- CP-element group 13: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Sample/word_access_start/$exit
      -- 
    ra_7555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2673_load_0_ack_0, ack => convTransposeD_CP_7276_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (12) 
      -- CP-element group 14: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2677_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Update/ptr_deref_2673_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Update/ptr_deref_2673_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Update/ptr_deref_2673_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Update/ptr_deref_2673_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2673_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2677_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2677_Sample/rr
      -- 
    ca_7566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2673_load_0_ack_1, ack => convTransposeD_CP_7276_elements(14)); -- 
    rr_7579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(14), ack => type_cast_2677_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2677_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2677_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2677_Sample/$exit
      -- 
    ra_7580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2677_inst_ack_0, ack => convTransposeD_CP_7276_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	33 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2677_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2677_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2677_update_completed_
      -- 
    ca_7585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2677_inst_ack_1, ack => convTransposeD_CP_7276_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Sample/word_access_start/word_0/ra
      -- 
    ra_7619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2689_load_0_ack_0, ack => convTransposeD_CP_7276_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	33 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Update/ptr_deref_2689_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Update/ptr_deref_2689_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Update/ptr_deref_2689_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2689_Update/ptr_deref_2689_Merge/$exit
      -- 
    ca_7630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2689_load_0_ack_1, ack => convTransposeD_CP_7276_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Sample/word_access_start/word_0/ra
      -- CP-element group 19: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Sample/word_access_start/word_0/$exit
      -- 
    ra_7652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2692_load_0_ack_0, ack => convTransposeD_CP_7276_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (12) 
      -- CP-element group 20: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Update/LOAD_padding_2692_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Update/LOAD_padding_2692_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2696_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Update/LOAD_padding_2692_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Update/LOAD_padding_2692_Merge/merge_ack
      -- CP-element group 20: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/LOAD_padding_2692_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2696_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2696_Sample/rr
      -- 
    ca_7663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2692_load_0_ack_1, ack => convTransposeD_CP_7276_elements(20)); -- 
    rr_7676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(20), ack => type_cast_2696_inst_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2696_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2696_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2696_Sample/$exit
      -- 
    ra_7677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2696_inst_ack_0, ack => convTransposeD_CP_7276_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	33 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2696_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2696_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2696_update_completed_
      -- 
    ca_7682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2696_inst_ack_1, ack => convTransposeD_CP_7276_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Sample/word_access_start/word_0/ra
      -- 
    ra_7716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2706_load_0_ack_0, ack => convTransposeD_CP_7276_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (12) 
      -- CP-element group 24: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Update/ptr_deref_2706_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Update/ptr_deref_2706_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Update/ptr_deref_2706_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2706_Update/ptr_deref_2706_Merge/merge_ack
      -- CP-element group 24: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2710_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2710_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2710_Sample/rr
      -- 
    ca_7727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2706_load_0_ack_1, ack => convTransposeD_CP_7276_elements(24)); -- 
    rr_7740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(24), ack => type_cast_2710_inst_req_0); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2710_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2710_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2710_Sample/ra
      -- 
    ra_7741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2710_inst_ack_0, ack => convTransposeD_CP_7276_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	33 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2710_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2710_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/type_cast_2710_Update/ca
      -- 
    ca_7746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2710_inst_ack_1, ack => convTransposeD_CP_7276_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Sample/word_access_start/word_0/ra
      -- 
    ra_7780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2722_load_0_ack_0, ack => convTransposeD_CP_7276_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	33 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Update/ptr_deref_2722_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Update/ptr_deref_2722_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Update/ptr_deref_2722_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2722_Update/ptr_deref_2722_Merge/merge_ack
      -- 
    ca_7791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2722_load_0_ack_1, ack => convTransposeD_CP_7276_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Sample/word_access_start/word_0/ra
      -- 
    ra_7830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2734_load_0_ack_0, ack => convTransposeD_CP_7276_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Update/ptr_deref_2734_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Update/ptr_deref_2734_Merge/$exit
      -- CP-element group 30: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Update/ptr_deref_2734_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2734_Update/ptr_deref_2734_Merge/merge_ack
      -- 
    ca_7841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2734_load_0_ack_1, ack => convTransposeD_CP_7276_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	2 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Sample/word_access_start/$exit
      -- CP-element group 31: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Sample/word_access_start/word_0/ra
      -- 
    ra_7880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2746_load_0_ack_0, ack => convTransposeD_CP_7276_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	2 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (9) 
      -- CP-element group 32: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Update/word_access_complete/$exit
      -- CP-element group 32: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Update/word_access_complete/word_0/ca
      -- CP-element group 32: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Update/ptr_deref_2746_Merge/$entry
      -- CP-element group 32: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Update/ptr_deref_2746_Merge/$exit
      -- CP-element group 32: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Update/ptr_deref_2746_Merge/merge_req
      -- CP-element group 32: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/ptr_deref_2746_Update/ptr_deref_2746_Merge/merge_ack
      -- 
    ca_7891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2746_load_0_ack_1, ack => convTransposeD_CP_7276_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  place  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: 	26 
    -- CP-element group 33: 	22 
    -- CP-element group 33: 	16 
    -- CP-element group 33: 	28 
    -- CP-element group 33: 	30 
    -- CP-element group 33: 	18 
    -- CP-element group 33: 	6 
    -- CP-element group 33: 	10 
    -- CP-element group 33: 	12 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	76 
    -- CP-element group 33: 	75 
    -- CP-element group 33: 	78 
    -- CP-element group 33: 	79 
    -- CP-element group 33:  members (20) 
      -- CP-element group 33: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747__exit__
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter
      -- CP-element group 33: 	 branch_block_stmt_2604/assign_stmt_2616_to_assign_stmt_2747/$exit
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/$entry
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2753/$entry
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2753/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2753/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2753/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2753/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2753/SplitProtocol/Update/cr
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/$entry
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/$entry
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Update/cr
      -- 
    rr_8325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(33), ack => type_cast_2753_inst_req_0); -- 
    cr_8330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(33), ack => type_cast_2753_inst_req_1); -- 
    rr_8348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(33), ack => type_cast_2759_inst_req_0); -- 
    cr_8353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(33), ack => type_cast_2759_inst_req_1); -- 
    convTransposeD_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(32) & convTransposeD_CP_7276_elements(26) & convTransposeD_CP_7276_elements(22) & convTransposeD_CP_7276_elements(16) & convTransposeD_CP_7276_elements(28) & convTransposeD_CP_7276_elements(30) & convTransposeD_CP_7276_elements(18) & convTransposeD_CP_7276_elements(6) & convTransposeD_CP_7276_elements(10) & convTransposeD_CP_7276_elements(12);
      gj_convTransposeD_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	92 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2766_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2766_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2766_Sample/ra
      -- 
    ra_7908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2766_inst_ack_0, ack => convTransposeD_CP_7276_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	92 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2766_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2766_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2766_Update/ca
      -- 
    ca_7913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2766_inst_ack_1, ack => convTransposeD_CP_7276_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	92 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2771_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2771_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2771_Sample/ra
      -- 
    ra_7922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2771_inst_ack_0, ack => convTransposeD_CP_7276_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	92 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2771_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2771_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2771_Update/ca
      -- 
    ca_7927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2771_inst_ack_1, ack => convTransposeD_CP_7276_elements(37)); -- 
    -- CP-element group 38:  join  transition  place  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	96 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874__exit__
      -- CP-element group 38: 	 branch_block_stmt_2604/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 38: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/$exit
      -- CP-element group 38: 	 branch_block_stmt_2604/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 38: 	 branch_block_stmt_2604/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2877/$entry
      -- CP-element group 38: 	 branch_block_stmt_2604/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/$entry
      -- 
    convTransposeD_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(35) & convTransposeD_CP_7276_elements(37);
      gj_convTransposeD_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	98 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2893_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2893_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2893_Sample/ra
      -- 
    ra_7939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2893_inst_ack_0, ack => convTransposeD_CP_7276_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	98 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	49 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (9) 
      -- CP-element group 40: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2893_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2893_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2893_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2923_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2923_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2923_Sample/rr
      -- CP-element group 40: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2954_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2954_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2954_Sample/rr
      -- 
    ca_7944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2893_inst_ack_1, ack => convTransposeD_CP_7276_elements(40)); -- 
    rr_8062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(40), ack => type_cast_2954_inst_req_0); -- 
    rr_7952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(40), ack => type_cast_2923_inst_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2923_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2923_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2923_Sample/ra
      -- 
    ra_7953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2923_inst_ack_0, ack => convTransposeD_CP_7276_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	98 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (16) 
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2923_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2923_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2923_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_index_resized_1
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_index_scaled_1
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_index_computed_1
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_index_resize_1/$entry
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_index_resize_1/$exit
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_index_resize_1/index_resize_req
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_index_resize_1/index_resize_ack
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_index_scale_1/$entry
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_index_scale_1/$exit
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_index_scale_1/scale_rename_req
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_index_scale_1/scale_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_final_index_sum_regn_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_final_index_sum_regn_Sample/req
      -- 
    ca_7958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2923_inst_ack_1, ack => convTransposeD_CP_7276_elements(42)); -- 
    req_7983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(42), ack => array_obj_ref_2929_index_offset_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	60 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_final_index_sum_regn_sample_complete
      -- CP-element group 43: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_final_index_sum_regn_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_final_index_sum_regn_Sample/ack
      -- 
    ack_7984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2929_index_offset_ack_0, ack => convTransposeD_CP_7276_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	98 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (11) 
      -- CP-element group 44: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2930_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_offset_calculated
      -- CP-element group 44: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_final_index_sum_regn_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_final_index_sum_regn_Update/ack
      -- CP-element group 44: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2930_request/$entry
      -- CP-element group 44: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2930_request/req
      -- 
    ack_7989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2929_index_offset_ack_1, ack => convTransposeD_CP_7276_elements(44)); -- 
    req_7998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(44), ack => addr_of_2930_final_reg_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2930_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2930_request/$exit
      -- CP-element group 45: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2930_request/ack
      -- 
    ack_7999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2930_final_reg_ack_0, ack => convTransposeD_CP_7276_elements(45)); -- 
    -- CP-element group 46:  join  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	98 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (24) 
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2930_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2930_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2930_complete/ack
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_base_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_word_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_root_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_base_address_resized
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_base_addr_resize/$entry
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_base_addr_resize/$exit
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_base_addr_resize/base_resize_req
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_base_addr_resize/base_resize_ack
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_base_plus_offset/$entry
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_base_plus_offset/$exit
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_base_plus_offset/sum_rename_req
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_base_plus_offset/sum_rename_ack
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_word_addrgen/$entry
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_word_addrgen/$exit
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_word_addrgen/root_register_req
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_word_addrgen/root_register_ack
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Sample/word_access_start/$entry
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Sample/word_access_start/word_0/$entry
      -- CP-element group 46: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Sample/word_access_start/word_0/rr
      -- 
    ack_8004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2930_final_reg_ack_1, ack => convTransposeD_CP_7276_elements(46)); -- 
    rr_8037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(46), ack => ptr_deref_2934_load_0_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (5) 
      -- CP-element group 47: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Sample/word_access_start/$exit
      -- CP-element group 47: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Sample/word_access_start/word_0/$exit
      -- CP-element group 47: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Sample/word_access_start/word_0/ra
      -- 
    ra_8038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2934_load_0_ack_0, ack => convTransposeD_CP_7276_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	98 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	55 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Update/word_access_complete/$exit
      -- CP-element group 48: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Update/word_access_complete/word_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Update/word_access_complete/word_0/ca
      -- CP-element group 48: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Update/ptr_deref_2934_Merge/$entry
      -- CP-element group 48: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Update/ptr_deref_2934_Merge/$exit
      -- CP-element group 48: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Update/ptr_deref_2934_Merge/merge_req
      -- CP-element group 48: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Update/ptr_deref_2934_Merge/merge_ack
      -- 
    ca_8049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2934_load_0_ack_1, ack => convTransposeD_CP_7276_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	40 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2954_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2954_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2954_Sample/ra
      -- 
    ra_8063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2954_inst_ack_0, ack => convTransposeD_CP_7276_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	98 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (16) 
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2954_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2954_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2954_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_index_resized_1
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_index_scaled_1
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_index_computed_1
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_index_resize_1/$entry
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_index_resize_1/$exit
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_index_resize_1/index_resize_req
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_index_resize_1/index_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_index_scale_1/$entry
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_index_scale_1/$exit
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_index_scale_1/scale_rename_req
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_index_scale_1/scale_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_final_index_sum_regn_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_final_index_sum_regn_Sample/req
      -- 
    ca_8068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2954_inst_ack_1, ack => convTransposeD_CP_7276_elements(50)); -- 
    req_8093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(50), ack => array_obj_ref_2960_index_offset_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	60 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_final_index_sum_regn_sample_complete
      -- CP-element group 51: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_final_index_sum_regn_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_final_index_sum_regn_Sample/ack
      -- 
    ack_8094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2960_index_offset_ack_0, ack => convTransposeD_CP_7276_elements(51)); -- 
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	98 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (11) 
      -- CP-element group 52: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2961_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_offset_calculated
      -- CP-element group 52: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_final_index_sum_regn_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_final_index_sum_regn_Update/ack
      -- CP-element group 52: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2961_request/$entry
      -- CP-element group 52: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2961_request/req
      -- 
    ack_8099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2960_index_offset_ack_1, ack => convTransposeD_CP_7276_elements(52)); -- 
    req_8108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(52), ack => addr_of_2961_final_reg_req_0); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2961_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2961_request/$exit
      -- CP-element group 53: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2961_request/ack
      -- 
    ack_8109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2961_final_reg_ack_0, ack => convTransposeD_CP_7276_elements(53)); -- 
    -- CP-element group 54:  fork  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	98 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (19) 
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2961_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2961_complete/$exit
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2961_complete/ack
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_base_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_word_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_root_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_base_address_resized
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_base_addr_resize/$entry
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_base_addr_resize/$exit
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_base_addr_resize/base_resize_req
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_base_addr_resize/base_resize_ack
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_base_plus_offset/$entry
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_base_plus_offset/$exit
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_base_plus_offset/sum_rename_req
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_base_plus_offset/sum_rename_ack
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_word_addrgen/$entry
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_word_addrgen/$exit
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_word_addrgen/root_register_req
      -- CP-element group 54: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_word_addrgen/root_register_ack
      -- 
    ack_8114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2961_final_reg_ack_1, ack => convTransposeD_CP_7276_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: 	48 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Sample/ptr_deref_2964_Split/$entry
      -- CP-element group 55: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Sample/ptr_deref_2964_Split/$exit
      -- CP-element group 55: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Sample/ptr_deref_2964_Split/split_req
      -- CP-element group 55: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Sample/ptr_deref_2964_Split/split_ack
      -- CP-element group 55: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Sample/word_access_start/word_0/rr
      -- 
    rr_8152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(55), ack => ptr_deref_2964_store_0_req_0); -- 
    convTransposeD_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(54) & convTransposeD_CP_7276_elements(48);
      gj_convTransposeD_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Sample/word_access_start/word_0/ra
      -- 
    ra_8153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2964_store_0_ack_0, ack => convTransposeD_CP_7276_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	98 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	60 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Update/word_access_complete/word_0/ca
      -- 
    ca_8164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2964_store_0_ack_1, ack => convTransposeD_CP_7276_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	98 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2970_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2970_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2970_Sample/ra
      -- 
    ra_8173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2970_inst_ack_0, ack => convTransposeD_CP_7276_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	98 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2970_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2970_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2970_Update/ca
      -- 
    ca_8178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2970_inst_ack_1, ack => convTransposeD_CP_7276_elements(59)); -- 
    -- CP-element group 60:  branch  join  transition  place  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: 	43 
    -- CP-element group 60: 	57 
    -- CP-element group 60: 	51 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (10) 
      -- CP-element group 60: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982__exit__
      -- CP-element group 60: 	 branch_block_stmt_2604/if_stmt_2983__entry__
      -- CP-element group 60: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/$exit
      -- CP-element group 60: 	 branch_block_stmt_2604/if_stmt_2983_dead_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_2604/if_stmt_2983_eval_test/$entry
      -- CP-element group 60: 	 branch_block_stmt_2604/if_stmt_2983_eval_test/$exit
      -- CP-element group 60: 	 branch_block_stmt_2604/if_stmt_2983_eval_test/branch_req
      -- CP-element group 60: 	 branch_block_stmt_2604/R_cmp_2984_place
      -- CP-element group 60: 	 branch_block_stmt_2604/if_stmt_2983_if_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_2604/if_stmt_2983_else_link/$entry
      -- 
    branch_req_8186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(60), ack => if_stmt_2983_branch_req_0); -- 
    convTransposeD_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(59) & convTransposeD_CP_7276_elements(43) & convTransposeD_CP_7276_elements(57) & convTransposeD_CP_7276_elements(51);
      gj_convTransposeD_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	93 
    -- CP-element group 61: 	94 
    -- CP-element group 61:  members (24) 
      -- CP-element group 61: 	 branch_block_stmt_2604/merge_stmt_2989__exit__
      -- CP-element group 61: 	 branch_block_stmt_2604/assign_stmt_2995__entry__
      -- CP-element group 61: 	 branch_block_stmt_2604/assign_stmt_2995__exit__
      -- CP-element group 61: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody
      -- CP-element group 61: 	 branch_block_stmt_2604/if_stmt_2983_if_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_2604/if_stmt_2983_if_link/if_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_2604/whilex_xbody_ifx_xthen
      -- CP-element group 61: 	 branch_block_stmt_2604/assign_stmt_2995/$entry
      -- CP-element group 61: 	 branch_block_stmt_2604/assign_stmt_2995/$exit
      -- CP-element group 61: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/$entry
      -- CP-element group 61: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/type_cast_2883/$entry
      -- CP-element group 61: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/type_cast_2883/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/type_cast_2883/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/type_cast_2883/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/type_cast_2883/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/type_cast_2883/SplitProtocol/Update/cr
      -- CP-element group 61: 	 branch_block_stmt_2604/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_2604/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 61: 	 branch_block_stmt_2604/merge_stmt_2989_PhiReqMerge
      -- CP-element group 61: 	 branch_block_stmt_2604/merge_stmt_2989_PhiAck/$entry
      -- CP-element group 61: 	 branch_block_stmt_2604/merge_stmt_2989_PhiAck/$exit
      -- CP-element group 61: 	 branch_block_stmt_2604/merge_stmt_2989_PhiAck/dummy
      -- 
    if_choice_transition_8191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2983_branch_ack_1, ack => convTransposeD_CP_7276_elements(61)); -- 
    rr_8429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(61), ack => type_cast_2883_inst_req_0); -- 
    cr_8434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(61), ack => type_cast_2883_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (18) 
      -- CP-element group 62: 	 branch_block_stmt_2604/merge_stmt_2997__exit__
      -- CP-element group 62: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013__entry__
      -- CP-element group 62: 	 branch_block_stmt_2604/if_stmt_2983_else_link/$exit
      -- CP-element group 62: 	 branch_block_stmt_2604/if_stmt_2983_else_link/else_choice_transition
      -- CP-element group 62: 	 branch_block_stmt_2604/whilex_xbody_ifx_xelse
      -- CP-element group 62: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/$entry
      -- CP-element group 62: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/type_cast_3007_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/type_cast_3007_update_start_
      -- CP-element group 62: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/type_cast_3007_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/type_cast_3007_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/type_cast_3007_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/type_cast_3007_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_2604/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 62: 	 branch_block_stmt_2604/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_2604/merge_stmt_2997_PhiReqMerge
      -- CP-element group 62: 	 branch_block_stmt_2604/merge_stmt_2997_PhiAck/$entry
      -- CP-element group 62: 	 branch_block_stmt_2604/merge_stmt_2997_PhiAck/$exit
      -- CP-element group 62: 	 branch_block_stmt_2604/merge_stmt_2997_PhiAck/dummy
      -- 
    else_choice_transition_8195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2983_branch_ack_0, ack => convTransposeD_CP_7276_elements(62)); -- 
    rr_8211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(62), ack => type_cast_3007_inst_req_0); -- 
    cr_8216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(62), ack => type_cast_3007_inst_req_1); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/type_cast_3007_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/type_cast_3007_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/type_cast_3007_Sample/ra
      -- 
    ra_8212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3007_inst_ack_0, ack => convTransposeD_CP_7276_elements(63)); -- 
    -- CP-element group 64:  branch  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (13) 
      -- CP-element group 64: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013__exit__
      -- CP-element group 64: 	 branch_block_stmt_2604/if_stmt_3014__entry__
      -- CP-element group 64: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/$exit
      -- CP-element group 64: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/type_cast_3007_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/type_cast_3007_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2604/assign_stmt_3003_to_assign_stmt_3013/type_cast_3007_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_2604/if_stmt_3014_dead_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_2604/if_stmt_3014_eval_test/$entry
      -- CP-element group 64: 	 branch_block_stmt_2604/if_stmt_3014_eval_test/$exit
      -- CP-element group 64: 	 branch_block_stmt_2604/if_stmt_3014_eval_test/branch_req
      -- CP-element group 64: 	 branch_block_stmt_2604/R_cmp81_3015_place
      -- CP-element group 64: 	 branch_block_stmt_2604/if_stmt_3014_if_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_2604/if_stmt_3014_else_link/$entry
      -- 
    ca_8217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3007_inst_ack_1, ack => convTransposeD_CP_7276_elements(64)); -- 
    branch_req_8225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(64), ack => if_stmt_3014_branch_req_0); -- 
    -- CP-element group 65:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (18) 
      -- CP-element group 65: 	 branch_block_stmt_2604/merge_stmt_3020__exit__
      -- CP-element group 65: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036__entry__
      -- CP-element group 65: 	 branch_block_stmt_2604/if_stmt_3014_if_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_2604/if_stmt_3014_if_link/if_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_2604/ifx_xelse_ifx_xthen83
      -- CP-element group 65: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/$entry
      -- CP-element group 65: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/type_cast_3035_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/type_cast_3035_update_start_
      -- CP-element group 65: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/type_cast_3035_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/type_cast_3035_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/type_cast_3035_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/type_cast_3035_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_2604/ifx_xelse_ifx_xthen83_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_2604/ifx_xelse_ifx_xthen83_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_2604/merge_stmt_3020_PhiReqMerge
      -- CP-element group 65: 	 branch_block_stmt_2604/merge_stmt_3020_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_2604/merge_stmt_3020_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_2604/merge_stmt_3020_PhiAck/dummy
      -- 
    if_choice_transition_8230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3014_branch_ack_1, ack => convTransposeD_CP_7276_elements(65)); -- 
    rr_8247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(65), ack => type_cast_3035_inst_req_0); -- 
    cr_8252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(65), ack => type_cast_3035_inst_req_1); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	99 
    -- CP-element group 66: 	100 
    -- CP-element group 66: 	102 
    -- CP-element group 66: 	103 
    -- CP-element group 66:  members (20) 
      -- CP-element group 66: 	 branch_block_stmt_2604/if_stmt_3014_else_link/$exit
      -- CP-element group 66: 	 branch_block_stmt_2604/if_stmt_3014_else_link/else_choice_transition
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/$entry
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3044/$entry
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3044/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3044/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3044/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3044/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3044/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/$entry
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3050/$entry
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3050/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3050/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3050/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3050/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3050/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3014_branch_ack_0, ack => convTransposeD_CP_7276_elements(66)); -- 
    rr_8503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(66), ack => type_cast_3044_inst_req_0); -- 
    cr_8508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(66), ack => type_cast_3044_inst_req_1); -- 
    rr_8526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(66), ack => type_cast_3050_inst_req_0); -- 
    cr_8531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(66), ack => type_cast_3050_inst_req_1); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/type_cast_3035_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/type_cast_3035_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/type_cast_3035_Sample/ra
      -- 
    ra_8248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3035_inst_ack_0, ack => convTransposeD_CP_7276_elements(67)); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	65 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	109 
    -- CP-element group 68: 	110 
    -- CP-element group 68: 	106 
    -- CP-element group 68: 	107 
    -- CP-element group 68:  members (23) 
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3048/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3048/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3042/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3042/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3042/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036__exit__
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3048/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3048/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3048/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3042/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3042/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3048/$entry
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/$entry
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3042/$entry
      -- CP-element group 68: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/$exit
      -- CP-element group 68: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/type_cast_3035_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/type_cast_3035_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_2604/assign_stmt_3026_to_assign_stmt_3036/type_cast_3035_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/$entry
      -- CP-element group 68: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/$entry
      -- 
    ca_8253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3035_inst_ack_1, ack => convTransposeD_CP_7276_elements(68)); -- 
    cr_8580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(68), ack => type_cast_3048_inst_req_1); -- 
    rr_8552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(68), ack => type_cast_3042_inst_req_0); -- 
    cr_8557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(68), ack => type_cast_3042_inst_req_1); -- 
    rr_8575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(68), ack => type_cast_3048_inst_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	116 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/type_cast_3055_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/type_cast_3055_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/type_cast_3055_Sample/ra
      -- 
    ra_8265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3055_inst_ack_0, ack => convTransposeD_CP_7276_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	116 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061__exit__
      -- CP-element group 70: 	 branch_block_stmt_2604/if_stmt_3062__entry__
      -- CP-element group 70: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/$exit
      -- CP-element group 70: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/type_cast_3055_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/type_cast_3055_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/type_cast_3055_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2604/if_stmt_3062_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2604/if_stmt_3062_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2604/if_stmt_3062_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2604/if_stmt_3062_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2604/R_cmp92_3063_place
      -- CP-element group 70: 	 branch_block_stmt_2604/if_stmt_3062_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2604/if_stmt_3062_else_link/$entry
      -- 
    ca_8270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3055_inst_ack_1, ack => convTransposeD_CP_7276_elements(70)); -- 
    branch_req_8278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(70), ack => if_stmt_3062_branch_req_0); -- 
    -- CP-element group 71:  merge  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2604/ifx_xend_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2604/ifx_xend_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2604/merge_stmt_3068_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2604/merge_stmt_3068_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2604/merge_stmt_3068_PhiAck/dummy
      -- CP-element group 71: 	 branch_block_stmt_2604/merge_stmt_3068__exit__
      -- CP-element group 71: 	 branch_block_stmt_2604/assign_stmt_3072__entry__
      -- CP-element group 71: 	 branch_block_stmt_2604/merge_stmt_3068_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2604/if_stmt_3062_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2604/if_stmt_3062_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2604/ifx_xend_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2604/assign_stmt_3072/$entry
      -- CP-element group 71: 	 branch_block_stmt_2604/assign_stmt_3072/WPIPE_Block3_done_3070_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2604/assign_stmt_3072/WPIPE_Block3_done_3070_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2604/assign_stmt_3072/WPIPE_Block3_done_3070_Sample/req
      -- 
    if_choice_transition_8283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3062_branch_ack_1, ack => convTransposeD_CP_7276_elements(71)); -- 
    req_8300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(71), ack => WPIPE_Block3_done_3070_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	82 
    -- CP-element group 72: 	83 
    -- CP-element group 72: 	85 
    -- CP-element group 72: 	86 
    -- CP-element group 72:  members (20) 
      -- CP-element group 72: 	 branch_block_stmt_2604/if_stmt_3062_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2604/if_stmt_3062_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/$entry
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2755/$entry
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2755/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2755/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2755/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2755/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2755/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/$entry
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2761/$entry
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2761/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2761/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2761/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2761/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2761/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3062_branch_ack_0, ack => convTransposeD_CP_7276_elements(72)); -- 
    rr_8374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(72), ack => type_cast_2755_inst_req_0); -- 
    cr_8379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(72), ack => type_cast_2755_inst_req_1); -- 
    rr_8397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(72), ack => type_cast_2761_inst_req_0); -- 
    cr_8402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(72), ack => type_cast_2761_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2604/assign_stmt_3072/WPIPE_Block3_done_3070_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2604/assign_stmt_3072/WPIPE_Block3_done_3070_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2604/assign_stmt_3072/WPIPE_Block3_done_3070_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2604/assign_stmt_3072/WPIPE_Block3_done_3070_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2604/assign_stmt_3072/WPIPE_Block3_done_3070_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2604/assign_stmt_3072/WPIPE_Block3_done_3070_Update/req
      -- 
    ack_8301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3070_inst_ack_0, ack => convTransposeD_CP_7276_elements(73)); -- 
    req_8305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(73), ack => WPIPE_Block3_done_3070_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2604/$exit
      -- CP-element group 74: 	 branch_block_stmt_2604/branch_block_stmt_2604__exit__
      -- CP-element group 74: 	 branch_block_stmt_2604/assign_stmt_3072__exit__
      -- CP-element group 74: 	 branch_block_stmt_2604/return__
      -- CP-element group 74: 	 branch_block_stmt_2604/merge_stmt_3074__exit__
      -- CP-element group 74: 	 branch_block_stmt_2604/merge_stmt_3074_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2604/merge_stmt_3074_PhiAck/dummy
      -- CP-element group 74: 	 branch_block_stmt_2604/merge_stmt_3074_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2604/merge_stmt_3074_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2604/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2604/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2604/assign_stmt_3072/$exit
      -- CP-element group 74: 	 branch_block_stmt_2604/assign_stmt_3072/WPIPE_Block3_done_3070_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2604/assign_stmt_3072/WPIPE_Block3_done_3070_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2604/assign_stmt_3072/WPIPE_Block3_done_3070_Update/ack
      -- 
    ack_8306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3070_inst_ack_1, ack => convTransposeD_CP_7276_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	33 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2753/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2753/SplitProtocol/Sample/ra
      -- 
    ra_8326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2753_inst_ack_0, ack => convTransposeD_CP_7276_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	33 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2753/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2753/SplitProtocol/Update/ca
      -- 
    ca_8331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2753_inst_ack_1, ack => convTransposeD_CP_7276_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/$exit
      -- CP-element group 77: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2753/$exit
      -- CP-element group 77: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2753/SplitProtocol/$exit
      -- CP-element group 77: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_req
      -- 
    phi_stmt_2750_req_8332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2750_req_8332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(77), ack => phi_stmt_2750_req_0); -- 
    convTransposeD_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(76) & convTransposeD_CP_7276_elements(75);
      gj_convTransposeD_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	33 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Sample/ra
      -- 
    ra_8349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2759_inst_ack_0, ack => convTransposeD_CP_7276_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	33 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Update/ca
      -- 
    ca_8354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2759_inst_ack_1, ack => convTransposeD_CP_7276_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/$exit
      -- CP-element group 80: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/$exit
      -- CP-element group 80: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_req
      -- 
    phi_stmt_2756_req_8355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2756_req_8355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(80), ack => phi_stmt_2756_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(78) & convTransposeD_CP_7276_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	89 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2604/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(77) & convTransposeD_CP_7276_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	72 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2755/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2755/SplitProtocol/Sample/ra
      -- 
    ra_8375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2755_inst_ack_0, ack => convTransposeD_CP_7276_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	72 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2755/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2755/SplitProtocol/Update/ca
      -- 
    ca_8380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2755_inst_ack_1, ack => convTransposeD_CP_7276_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	88 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/$exit
      -- CP-element group 84: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2755/$exit
      -- CP-element group 84: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_sources/type_cast_2755/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2750/phi_stmt_2750_req
      -- 
    phi_stmt_2750_req_8381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2750_req_8381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(84), ack => phi_stmt_2750_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(82) & convTransposeD_CP_7276_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	72 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2761/SplitProtocol/Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2761/SplitProtocol/Sample/ra
      -- 
    ra_8398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2761_inst_ack_0, ack => convTransposeD_CP_7276_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	72 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2761/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2761/SplitProtocol/Update/ca
      -- 
    ca_8403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2761_inst_ack_1, ack => convTransposeD_CP_7276_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/$exit
      -- CP-element group 87: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2761/$exit
      -- CP-element group 87: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2761/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2756/phi_stmt_2756_req
      -- 
    phi_stmt_2756_req_8404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2756_req_8404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(87), ack => phi_stmt_2756_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(85) & convTransposeD_CP_7276_elements(86);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  join  transition  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	84 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2604/ifx_xend_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(84) & convTransposeD_CP_7276_elements(87);
      gj_convTransposeD_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  merge  fork  transition  place  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	81 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2604/merge_stmt_2749_PhiReqMerge
      -- CP-element group 89: 	 branch_block_stmt_2604/merge_stmt_2749_PhiAck/$entry
      -- 
    convTransposeD_CP_7276_elements(89) <= OrReduce(convTransposeD_CP_7276_elements(81) & convTransposeD_CP_7276_elements(88));
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_2604/merge_stmt_2749_PhiAck/phi_stmt_2750_ack
      -- 
    phi_stmt_2750_ack_8409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2750_ack_0, ack => convTransposeD_CP_7276_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_2604/merge_stmt_2749_PhiAck/phi_stmt_2756_ack
      -- 
    phi_stmt_2756_ack_8410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2756_ack_0, ack => convTransposeD_CP_7276_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  place  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	35 
    -- CP-element group 92: 	36 
    -- CP-element group 92: 	37 
    -- CP-element group 92: 	34 
    -- CP-element group 92:  members (16) 
      -- CP-element group 92: 	 branch_block_stmt_2604/merge_stmt_2749__exit__
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874__entry__
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/$entry
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2766_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2766_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2766_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2766_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2766_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2766_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2771_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2771_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2771_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2771_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2771_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2604/assign_stmt_2767_to_assign_stmt_2874/type_cast_2771_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2604/merge_stmt_2749_PhiAck/$exit
      -- 
    rr_7907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(92), ack => type_cast_2766_inst_req_0); -- 
    cr_7912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(92), ack => type_cast_2766_inst_req_1); -- 
    rr_7921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(92), ack => type_cast_2771_inst_req_0); -- 
    cr_7926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(92), ack => type_cast_2771_inst_req_1); -- 
    convTransposeD_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(90) & convTransposeD_CP_7276_elements(91);
      gj_convTransposeD_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	61 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/type_cast_2883/SplitProtocol/Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/type_cast_2883/SplitProtocol/Sample/ra
      -- 
    ra_8430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2883_inst_ack_0, ack => convTransposeD_CP_7276_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	61 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/type_cast_2883/SplitProtocol/Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/type_cast_2883/SplitProtocol/Update/ca
      -- 
    ca_8435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2883_inst_ack_1, ack => convTransposeD_CP_7276_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 95: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/$exit
      -- CP-element group 95: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/type_cast_2883/$exit
      -- CP-element group 95: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/type_cast_2883/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_2604/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_req
      -- 
    phi_stmt_2877_req_8436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2877_req_8436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(95), ack => phi_stmt_2877_req_1); -- 
    convTransposeD_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(93) & convTransposeD_CP_7276_elements(94);
      gj_convTransposeD_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  transition  output  delay-element  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	38 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_2604/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 96: 	 branch_block_stmt_2604/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2877/$exit
      -- CP-element group 96: 	 branch_block_stmt_2604/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/$exit
      -- CP-element group 96: 	 branch_block_stmt_2604/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_sources/type_cast_2881_konst_delay_trans
      -- CP-element group 96: 	 branch_block_stmt_2604/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2877/phi_stmt_2877_req
      -- 
    phi_stmt_2877_req_8447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2877_req_8447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(96), ack => phi_stmt_2877_req_0); -- 
    -- Element group convTransposeD_CP_7276_elements(96) is a control-delay.
    cp_element_96_delay: control_delay_element  generic map(name => " 96_delay", delay_value => 1)  port map(req => convTransposeD_CP_7276_elements(38), ack => convTransposeD_CP_7276_elements(96), clk => clk, reset =>reset);
    -- CP-element group 97:  merge  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_2604/merge_stmt_2876_PhiReqMerge
      -- CP-element group 97: 	 branch_block_stmt_2604/merge_stmt_2876_PhiAck/$entry
      -- 
    convTransposeD_CP_7276_elements(97) <= OrReduce(convTransposeD_CP_7276_elements(95) & convTransposeD_CP_7276_elements(96));
    -- CP-element group 98:  fork  transition  place  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	50 
    -- CP-element group 98: 	59 
    -- CP-element group 98: 	54 
    -- CP-element group 98: 	40 
    -- CP-element group 98: 	46 
    -- CP-element group 98: 	44 
    -- CP-element group 98: 	57 
    -- CP-element group 98: 	48 
    -- CP-element group 98: 	42 
    -- CP-element group 98: 	39 
    -- CP-element group 98: 	58 
    -- CP-element group 98: 	52 
    -- CP-element group 98:  members (45) 
      -- CP-element group 98: 	 branch_block_stmt_2604/merge_stmt_2876__exit__
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982__entry__
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2893_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2893_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2893_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2893_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2893_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2893_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2923_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2923_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2923_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2930_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_final_index_sum_regn_update_start
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_final_index_sum_regn_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2929_final_index_sum_regn_Update/req
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2930_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2930_complete/req
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Update/word_access_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Update/word_access_complete/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2934_Update/word_access_complete/word_0/cr
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2954_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2954_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2954_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2961_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_final_index_sum_regn_update_start
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_final_index_sum_regn_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/array_obj_ref_2960_final_index_sum_regn_Update/req
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2961_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/addr_of_2961_complete/req
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Update/word_access_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Update/word_access_complete/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/ptr_deref_2964_Update/word_access_complete/word_0/cr
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2970_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2970_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2970_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2970_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2970_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2604/assign_stmt_2890_to_assign_stmt_2982/type_cast_2970_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2604/merge_stmt_2876_PhiAck/$exit
      -- CP-element group 98: 	 branch_block_stmt_2604/merge_stmt_2876_PhiAck/phi_stmt_2877_ack
      -- 
    phi_stmt_2877_ack_8452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2877_ack_0, ack => convTransposeD_CP_7276_elements(98)); -- 
    rr_7938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(98), ack => type_cast_2893_inst_req_0); -- 
    cr_7943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(98), ack => type_cast_2893_inst_req_1); -- 
    cr_7957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(98), ack => type_cast_2923_inst_req_1); -- 
    req_7988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(98), ack => array_obj_ref_2929_index_offset_req_1); -- 
    req_8003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(98), ack => addr_of_2930_final_reg_req_1); -- 
    cr_8048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(98), ack => ptr_deref_2934_load_0_req_1); -- 
    cr_8067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(98), ack => type_cast_2954_inst_req_1); -- 
    req_8098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(98), ack => array_obj_ref_2960_index_offset_req_1); -- 
    req_8113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(98), ack => addr_of_2961_final_reg_req_1); -- 
    cr_8163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(98), ack => ptr_deref_2964_store_0_req_1); -- 
    rr_8172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(98), ack => type_cast_2970_inst_req_0); -- 
    cr_8177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(98), ack => type_cast_2970_inst_req_1); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	66 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3044/SplitProtocol/Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3044/SplitProtocol/Sample/ra
      -- 
    ra_8504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3044_inst_ack_0, ack => convTransposeD_CP_7276_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	66 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3044/SplitProtocol/Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3044/SplitProtocol/Update/ca
      -- 
    ca_8509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3044_inst_ack_1, ack => convTransposeD_CP_7276_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	105 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/$exit
      -- CP-element group 101: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3044/$exit
      -- CP-element group 101: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3044/SplitProtocol/$exit
      -- CP-element group 101: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_req
      -- 
    phi_stmt_3039_req_8510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3039_req_8510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(101), ack => phi_stmt_3039_req_1); -- 
    convTransposeD_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(99) & convTransposeD_CP_7276_elements(100);
      gj_convTransposeD_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	66 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3050/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3050/SplitProtocol/Sample/ra
      -- 
    ra_8527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3050_inst_ack_0, ack => convTransposeD_CP_7276_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	66 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3050/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3050/SplitProtocol/Update/ca
      -- 
    ca_8532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3050_inst_ack_1, ack => convTransposeD_CP_7276_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/$exit
      -- CP-element group 104: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3050/$exit
      -- CP-element group 104: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3050/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_req
      -- 
    phi_stmt_3045_req_8533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3045_req_8533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(104), ack => phi_stmt_3045_req_1); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(102) & convTransposeD_CP_7276_elements(103);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	101 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	113 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_2604/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(101) & convTransposeD_CP_7276_elements(104);
      gj_convTransposeD_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	68 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3042/SplitProtocol/Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3042/SplitProtocol/Sample/$exit
      -- 
    ra_8553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3042_inst_ack_0, ack => convTransposeD_CP_7276_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	68 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3042/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3042/SplitProtocol/Update/ca
      -- 
    ca_8558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3042_inst_ack_1, ack => convTransposeD_CP_7276_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_req
      -- CP-element group 108: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3042/$exit
      -- CP-element group 108: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/type_cast_3042/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/$exit
      -- CP-element group 108: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3039/phi_stmt_3039_sources/$exit
      -- 
    phi_stmt_3039_req_8559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3039_req_8559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(108), ack => phi_stmt_3039_req_0); -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(106) & convTransposeD_CP_7276_elements(107);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	68 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3048/SplitProtocol/Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3048/SplitProtocol/Sample/$exit
      -- 
    ra_8576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3048_inst_ack_0, ack => convTransposeD_CP_7276_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	68 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3048/SplitProtocol/Update/ca
      -- CP-element group 110: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3048/SplitProtocol/Update/$exit
      -- 
    ca_8581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3048_inst_ack_1, ack => convTransposeD_CP_7276_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_req
      -- CP-element group 111: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3048/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/type_cast_3048/$exit
      -- CP-element group 111: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/phi_stmt_3045_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3045/$exit
      -- 
    phi_stmt_3045_req_8582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3045_req_8582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(111), ack => phi_stmt_3045_req_0); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(109) & convTransposeD_CP_7276_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: 	108 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2604/ifx_xthen83_ifx_xend_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(111) & convTransposeD_CP_7276_elements(108);
      gj_convTransposeD_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  merge  fork  transition  place  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	105 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2604/merge_stmt_3038_PhiAck/$entry
      -- CP-element group 113: 	 branch_block_stmt_2604/merge_stmt_3038_PhiReqMerge
      -- 
    convTransposeD_CP_7276_elements(113) <= OrReduce(convTransposeD_CP_7276_elements(105) & convTransposeD_CP_7276_elements(112));
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_2604/merge_stmt_3038_PhiAck/phi_stmt_3039_ack
      -- 
    phi_stmt_3039_ack_8587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3039_ack_0, ack => convTransposeD_CP_7276_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_2604/merge_stmt_3038_PhiAck/phi_stmt_3045_ack
      -- 
    phi_stmt_3045_ack_8588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3045_ack_0, ack => convTransposeD_CP_7276_elements(115)); -- 
    -- CP-element group 116:  join  fork  transition  place  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: 	70 
    -- CP-element group 116:  members (10) 
      -- CP-element group 116: 	 branch_block_stmt_2604/merge_stmt_3038_PhiAck/$exit
      -- CP-element group 116: 	 branch_block_stmt_2604/merge_stmt_3038__exit__
      -- CP-element group 116: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061__entry__
      -- CP-element group 116: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/$entry
      -- CP-element group 116: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/type_cast_3055_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/type_cast_3055_update_start_
      -- CP-element group 116: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/type_cast_3055_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/type_cast_3055_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/type_cast_3055_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_2604/assign_stmt_3056_to_assign_stmt_3061/type_cast_3055_Update/cr
      -- 
    rr_8264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(116), ack => type_cast_3055_inst_req_0); -- 
    cr_8269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7276_elements(116), ack => type_cast_3055_inst_req_1); -- 
    convTransposeD_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7276_elements(114) & convTransposeD_CP_7276_elements(115);
      gj_convTransposeD_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7276_elements(116), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2836_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2857_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2917_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2948_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_2692_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2692_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom65_2959_resized : std_logic_vector(13 downto 0);
    signal R_idxprom65_2959_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2928_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2928_scaled : std_logic_vector(13 downto 0);
    signal add21_2899 : std_logic_vector(31 downto 0);
    signal add29_2797 : std_logic_vector(31 downto 0);
    signal add40_2812 : std_logic_vector(31 downto 0);
    signal add55_2869 : std_logic_vector(31 downto 0);
    signal add57_2904 : std_logic_vector(31 downto 0);
    signal add70_2977 : std_logic_vector(31 downto 0);
    signal add_2782 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2929_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2929_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2929_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2929_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2929_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2929_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2960_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2960_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2960_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2960_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2960_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2960_root_address : std_logic_vector(13 downto 0);
    signal arrayidx66_2962 : std_logic_vector(31 downto 0);
    signal arrayidx_2931 : std_logic_vector(31 downto 0);
    signal call_2607 : std_logic_vector(15 downto 0);
    signal cmp81_3013 : std_logic_vector(0 downto 0);
    signal cmp92_3061 : std_logic_vector(0 downto 0);
    signal cmp_2982 : std_logic_vector(0 downto 0);
    signal conv13105_2894 : std_logic_vector(31 downto 0);
    signal conv16_2767 : std_logic_vector(31 downto 0);
    signal conv19_2772 : std_logic_vector(31 downto 0);
    signal conv26_2678 : std_logic_vector(31 downto 0);
    signal conv31_2697 : std_logic_vector(31 downto 0);
    signal conv37_2711 : std_logic_vector(31 downto 0);
    signal conv4_2652 : std_logic_vector(15 downto 0);
    signal conv50_2838 : std_logic_vector(31 downto 0);
    signal conv53_2859 : std_logic_vector(31 downto 0);
    signal conv69_2971 : std_logic_vector(31 downto 0);
    signal conv79_3008 : std_logic_vector(31 downto 0);
    signal conv88_3036 : std_logic_vector(15 downto 0);
    signal conv90_3056 : std_logic_vector(31 downto 0);
    signal conv_2630 : std_logic_vector(15 downto 0);
    signal div3_2648 : std_logic_vector(31 downto 0);
    signal div87_3032 : std_logic_vector(31 downto 0);
    signal div_2626 : std_logic_vector(31 downto 0);
    signal iNsTr_10_2743 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2616 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2638 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2660 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2670 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2686 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2703 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2719 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2731 : std_logic_vector(31 downto 0);
    signal idxprom65_2955 : std_logic_vector(63 downto 0);
    signal idxprom_2924 : std_logic_vector(63 downto 0);
    signal inc85_3026 : std_logic_vector(15 downto 0);
    signal inc_3003 : std_logic_vector(15 downto 0);
    signal indvar_2877 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2995 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_3045 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2756 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2750 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_3039 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2890 : std_logic_vector(15 downto 0);
    signal mul20_2787 : std_logic_vector(31 downto 0);
    signal mul27_2792 : std_logic_vector(31 downto 0);
    signal mul38_2807 : std_logic_vector(31 downto 0);
    signal mul54_2864 : std_logic_vector(31 downto 0);
    signal mul56_2874 : std_logic_vector(31 downto 0);
    signal mul_2777 : std_logic_vector(31 downto 0);
    signal ptr_deref_2619_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2619_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2619_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2619_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2619_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2641_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2641_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2641_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2641_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2641_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2663_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2663_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2663_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2663_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2663_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2673_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2673_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2673_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2673_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2673_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2689_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2689_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2689_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2689_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2689_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2706_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2706_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2706_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2706_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2706_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2722_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2722_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2722_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2722_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2722_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2734_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2734_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2734_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2734_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2734_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2746_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2746_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2746_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2746_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2746_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2934_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2934_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2934_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2934_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2934_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2964_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2964_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2964_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2964_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2964_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2964_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext106_2850 : std_logic_vector(31 downto 0);
    signal sext108_2910 : std_logic_vector(31 downto 0);
    signal sext109_2941 : std_logic_vector(31 downto 0);
    signal sext_2829 : std_logic_vector(31 downto 0);
    signal shr64_2950 : std_logic_vector(31 downto 0);
    signal shr_2919 : std_logic_vector(31 downto 0);
    signal sub32_2844 : std_logic_vector(31 downto 0);
    signal sub43_2817 : std_logic_vector(31 downto 0);
    signal sub44_2823 : std_logic_vector(31 downto 0);
    signal sub_2802 : std_logic_vector(31 downto 0);
    signal tmp14_2664 : std_logic_vector(31 downto 0);
    signal tmp25_2674 : std_logic_vector(15 downto 0);
    signal tmp28_2690 : std_logic_vector(31 downto 0);
    signal tmp2_2642 : std_logic_vector(31 downto 0);
    signal tmp30_2693 : std_logic_vector(15 downto 0);
    signal tmp36_2707 : std_logic_vector(15 downto 0);
    signal tmp39_2723 : std_logic_vector(31 downto 0);
    signal tmp48_2735 : std_logic_vector(31 downto 0);
    signal tmp51_2747 : std_logic_vector(31 downto 0);
    signal tmp61_2935 : std_logic_vector(63 downto 0);
    signal tmp_2620 : std_logic_vector(31 downto 0);
    signal type_cast_2624_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2646_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2753_wire : std_logic_vector(15 downto 0);
    signal type_cast_2755_wire : std_logic_vector(15 downto 0);
    signal type_cast_2759_wire : std_logic_vector(15 downto 0);
    signal type_cast_2761_wire : std_logic_vector(15 downto 0);
    signal type_cast_2765_wire : std_logic_vector(31 downto 0);
    signal type_cast_2770_wire : std_logic_vector(31 downto 0);
    signal type_cast_2821_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2827_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2832_wire : std_logic_vector(31 downto 0);
    signal type_cast_2835_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2842_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2848_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2853_wire : std_logic_vector(31 downto 0);
    signal type_cast_2856_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2881_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2883_wire : std_logic_vector(15 downto 0);
    signal type_cast_2888_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2908_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2913_wire : std_logic_vector(31 downto 0);
    signal type_cast_2916_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2922_wire : std_logic_vector(63 downto 0);
    signal type_cast_2939_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2944_wire : std_logic_vector(31 downto 0);
    signal type_cast_2947_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2953_wire : std_logic_vector(63 downto 0);
    signal type_cast_2969_wire : std_logic_vector(31 downto 0);
    signal type_cast_2975_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2993_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3001_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3006_wire : std_logic_vector(31 downto 0);
    signal type_cast_3024_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3030_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3042_wire : std_logic_vector(15 downto 0);
    signal type_cast_3044_wire : std_logic_vector(15 downto 0);
    signal type_cast_3048_wire : std_logic_vector(15 downto 0);
    signal type_cast_3050_wire : std_logic_vector(15 downto 0);
    signal type_cast_3054_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_2692_word_address_0 <= "0";
    array_obj_ref_2929_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2929_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2929_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2929_resized_base_address <= "00000000000000";
    array_obj_ref_2960_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2960_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2960_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2960_resized_base_address <= "00000000000000";
    iNsTr_10_2743 <= "00000000000000000000000000000011";
    iNsTr_2_2616 <= "00000000000000000000000000000010";
    iNsTr_3_2638 <= "00000000000000000000000000000011";
    iNsTr_4_2660 <= "00000000000000000000000000000100";
    iNsTr_5_2670 <= "00000000000000000000000000000000";
    iNsTr_6_2686 <= "00000000000000000000000000000011";
    iNsTr_7_2703 <= "00000000000000000000000000000001";
    iNsTr_8_2719 <= "00000000000000000000000000000100";
    iNsTr_9_2731 <= "00000000000000000000000000000100";
    ptr_deref_2619_word_offset_0 <= "0000000";
    ptr_deref_2641_word_offset_0 <= "0000000";
    ptr_deref_2663_word_offset_0 <= "0000000";
    ptr_deref_2673_word_offset_0 <= "0";
    ptr_deref_2689_word_offset_0 <= "0000000";
    ptr_deref_2706_word_offset_0 <= "0";
    ptr_deref_2722_word_offset_0 <= "0000000";
    ptr_deref_2734_word_offset_0 <= "0000000";
    ptr_deref_2746_word_offset_0 <= "0000000";
    ptr_deref_2934_word_offset_0 <= "00000000000000";
    ptr_deref_2964_word_offset_0 <= "00000000000000";
    type_cast_2624_wire_constant <= "00000000000000000000000000000001";
    type_cast_2646_wire_constant <= "00000000000000000000000000000001";
    type_cast_2821_wire_constant <= "00000000000000000000000000010000";
    type_cast_2827_wire_constant <= "11111111111111110000000000000000";
    type_cast_2835_wire_constant <= "00000000000000000000000000010000";
    type_cast_2842_wire_constant <= "00000000000000000000000000010000";
    type_cast_2848_wire_constant <= "11111111111111110000000000000000";
    type_cast_2856_wire_constant <= "00000000000000000000000000010000";
    type_cast_2881_wire_constant <= "0000000000000000";
    type_cast_2888_wire_constant <= "0000000000000100";
    type_cast_2908_wire_constant <= "00000000000000000000000000010000";
    type_cast_2916_wire_constant <= "00000000000000000000000000010010";
    type_cast_2939_wire_constant <= "00000000000000000000000000010000";
    type_cast_2947_wire_constant <= "00000000000000000000000000010010";
    type_cast_2975_wire_constant <= "00000000000000000000000000000100";
    type_cast_2993_wire_constant <= "0000000000000001";
    type_cast_3001_wire_constant <= "0000000000000001";
    type_cast_3024_wire_constant <= "0000000000000001";
    type_cast_3030_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_2750: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2753_wire & type_cast_2755_wire;
      req <= phi_stmt_2750_req_0 & phi_stmt_2750_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2750",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2750_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2750,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2750
    phi_stmt_2756: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2759_wire & type_cast_2761_wire;
      req <= phi_stmt_2756_req_0 & phi_stmt_2756_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2756",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2756_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2756,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2756
    phi_stmt_2877: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2881_wire_constant & type_cast_2883_wire;
      req <= phi_stmt_2877_req_0 & phi_stmt_2877_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2877",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2877_ack_0,
          idata => idata,
          odata => indvar_2877,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2877
    phi_stmt_3039: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3042_wire & type_cast_3044_wire;
      req <= phi_stmt_3039_req_0 & phi_stmt_3039_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3039",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3039_ack_0,
          idata => idata,
          odata => input_dim1x_x2_3039,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3039
    phi_stmt_3045: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3048_wire & type_cast_3050_wire;
      req <= phi_stmt_3045_req_0 & phi_stmt_3045_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3045",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3045_ack_0,
          idata => idata,
          odata => input_dim0x_x0_3045,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3045
    addr_of_2930_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2930_final_reg_req_0;
      addr_of_2930_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2930_final_reg_req_1;
      addr_of_2930_final_reg_ack_1<= rack(0);
      addr_of_2930_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2930_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2929_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2931,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2961_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2961_final_reg_req_0;
      addr_of_2961_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2961_final_reg_req_1;
      addr_of_2961_final_reg_ack_1<= rack(0);
      addr_of_2961_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2961_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2960_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx66_2962,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2629_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2629_inst_req_0;
      type_cast_2629_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2629_inst_req_1;
      type_cast_2629_inst_ack_1<= rack(0);
      type_cast_2629_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2629_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2630,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2651_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2651_inst_req_0;
      type_cast_2651_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2651_inst_req_1;
      type_cast_2651_inst_ack_1<= rack(0);
      type_cast_2651_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2651_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div3_2648,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_2652,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2677_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2677_inst_req_0;
      type_cast_2677_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2677_inst_req_1;
      type_cast_2677_inst_ack_1<= rack(0);
      type_cast_2677_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2677_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp25_2674,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_2678,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2696_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2696_inst_req_0;
      type_cast_2696_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2696_inst_req_1;
      type_cast_2696_inst_ack_1<= rack(0);
      type_cast_2696_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2696_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp30_2693,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_2697,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2710_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2710_inst_req_0;
      type_cast_2710_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2710_inst_req_1;
      type_cast_2710_inst_ack_1<= rack(0);
      type_cast_2710_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2710_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp36_2707,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv37_2711,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2753_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2753_inst_req_0;
      type_cast_2753_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2753_inst_req_1;
      type_cast_2753_inst_ack_1<= rack(0);
      type_cast_2753_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2753_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_2652,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2753_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2755_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2755_inst_req_0;
      type_cast_2755_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2755_inst_req_1;
      type_cast_2755_inst_ack_1<= rack(0);
      type_cast_2755_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2755_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_3039,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2755_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2759_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2759_inst_req_0;
      type_cast_2759_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2759_inst_req_1;
      type_cast_2759_inst_ack_1<= rack(0);
      type_cast_2759_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2759_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_2630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2759_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2761_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2761_inst_req_0;
      type_cast_2761_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2761_inst_req_1;
      type_cast_2761_inst_ack_1<= rack(0);
      type_cast_2761_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2761_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_3045,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2761_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2766_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2766_inst_req_0;
      type_cast_2766_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2766_inst_req_1;
      type_cast_2766_inst_ack_1<= rack(0);
      type_cast_2766_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2766_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2765_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_2767,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2771_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2771_inst_req_0;
      type_cast_2771_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2771_inst_req_1;
      type_cast_2771_inst_ack_1<= rack(0);
      type_cast_2771_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2771_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2770_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_2772,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2832_inst
    process(sext_2829) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2829(31 downto 0);
      type_cast_2832_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2837_inst
    process(ASHR_i32_i32_2836_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2836_wire(31 downto 0);
      conv50_2838 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2853_inst
    process(sext106_2850) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext106_2850(31 downto 0);
      type_cast_2853_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2858_inst
    process(ASHR_i32_i32_2857_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2857_wire(31 downto 0);
      conv53_2859 <= tmp_var; -- 
    end process;
    type_cast_2883_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2883_inst_req_0;
      type_cast_2883_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2883_inst_req_1;
      type_cast_2883_inst_ack_1<= rack(0);
      type_cast_2883_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2883_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2995,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2883_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2893_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2893_inst_req_0;
      type_cast_2893_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2893_inst_req_1;
      type_cast_2893_inst_ack_1<= rack(0);
      type_cast_2893_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2893_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2890,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13105_2894,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2913_inst
    process(sext108_2910) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext108_2910(31 downto 0);
      type_cast_2913_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2918_inst
    process(ASHR_i32_i32_2917_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2917_wire(31 downto 0);
      shr_2919 <= tmp_var; -- 
    end process;
    type_cast_2923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2923_inst_req_0;
      type_cast_2923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2923_inst_req_1;
      type_cast_2923_inst_ack_1<= rack(0);
      type_cast_2923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2922_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2924,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2944_inst
    process(sext109_2941) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext109_2941(31 downto 0);
      type_cast_2944_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2949_inst
    process(ASHR_i32_i32_2948_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2948_wire(31 downto 0);
      shr64_2950 <= tmp_var; -- 
    end process;
    type_cast_2954_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2954_inst_req_0;
      type_cast_2954_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2954_inst_req_1;
      type_cast_2954_inst_ack_1<= rack(0);
      type_cast_2954_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2954_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2953_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom65_2955,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2970_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2970_inst_req_0;
      type_cast_2970_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2970_inst_req_1;
      type_cast_2970_inst_ack_1<= rack(0);
      type_cast_2970_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2970_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2969_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_2971,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3007_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3007_inst_req_0;
      type_cast_3007_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3007_inst_req_1;
      type_cast_3007_inst_ack_1<= rack(0);
      type_cast_3007_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3007_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3006_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_3008,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3035_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3035_inst_req_0;
      type_cast_3035_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3035_inst_req_1;
      type_cast_3035_inst_ack_1<= rack(0);
      type_cast_3035_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3035_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div87_3032,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv88_3036,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3042_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3042_inst_req_0;
      type_cast_3042_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3042_inst_req_1;
      type_cast_3042_inst_ack_1<= rack(0);
      type_cast_3042_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3042_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv88_3036,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3042_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3044_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3044_inst_req_0;
      type_cast_3044_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3044_inst_req_1;
      type_cast_3044_inst_ack_1<= rack(0);
      type_cast_3044_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3044_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_3003,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3044_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3048_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3048_inst_req_0;
      type_cast_3048_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3048_inst_req_1;
      type_cast_3048_inst_ack_1<= rack(0);
      type_cast_3048_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3048_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc85_3026,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3048_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3050_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3050_inst_req_0;
      type_cast_3050_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3050_inst_req_1;
      type_cast_3050_inst_ack_1<= rack(0);
      type_cast_3050_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3050_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2x_xph_2756,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3050_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3055_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3055_inst_req_0;
      type_cast_3055_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3055_inst_req_1;
      type_cast_3055_inst_ack_1<= rack(0);
      type_cast_3055_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3055_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3054_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_3056,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2692_gather_scatter
    process(LOAD_padding_2692_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2692_data_0;
      ov(15 downto 0) := iv;
      tmp30_2693 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2929_index_1_rename
    process(R_idxprom_2928_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2928_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2928_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2929_index_1_resize
    process(idxprom_2924) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2924;
      ov := iv(13 downto 0);
      R_idxprom_2928_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2929_root_address_inst
    process(array_obj_ref_2929_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2929_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2929_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2960_index_1_rename
    process(R_idxprom65_2959_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom65_2959_resized;
      ov(13 downto 0) := iv;
      R_idxprom65_2959_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2960_index_1_resize
    process(idxprom65_2955) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom65_2955;
      ov := iv(13 downto 0);
      R_idxprom65_2959_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2960_root_address_inst
    process(array_obj_ref_2960_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2960_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2960_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2619_addr_0
    process(ptr_deref_2619_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2619_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2619_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2619_base_resize
    process(iNsTr_2_2616) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2616;
      ov := iv(6 downto 0);
      ptr_deref_2619_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2619_gather_scatter
    process(ptr_deref_2619_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2619_data_0;
      ov(31 downto 0) := iv;
      tmp_2620 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2619_root_address_inst
    process(ptr_deref_2619_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2619_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2619_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2641_addr_0
    process(ptr_deref_2641_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2641_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2641_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2641_base_resize
    process(iNsTr_3_2638) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2638;
      ov := iv(6 downto 0);
      ptr_deref_2641_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2641_gather_scatter
    process(ptr_deref_2641_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2641_data_0;
      ov(31 downto 0) := iv;
      tmp2_2642 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2641_root_address_inst
    process(ptr_deref_2641_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2641_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2641_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2663_addr_0
    process(ptr_deref_2663_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2663_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2663_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2663_base_resize
    process(iNsTr_4_2660) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2660;
      ov := iv(6 downto 0);
      ptr_deref_2663_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2663_gather_scatter
    process(ptr_deref_2663_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2663_data_0;
      ov(31 downto 0) := iv;
      tmp14_2664 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2663_root_address_inst
    process(ptr_deref_2663_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2663_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2663_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2673_addr_0
    process(ptr_deref_2673_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2673_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2673_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2673_base_resize
    process(iNsTr_5_2670) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2670;
      ov := iv(0 downto 0);
      ptr_deref_2673_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2673_gather_scatter
    process(ptr_deref_2673_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2673_data_0;
      ov(15 downto 0) := iv;
      tmp25_2674 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2673_root_address_inst
    process(ptr_deref_2673_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2673_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2673_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2689_addr_0
    process(ptr_deref_2689_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2689_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2689_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2689_base_resize
    process(iNsTr_6_2686) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2686;
      ov := iv(6 downto 0);
      ptr_deref_2689_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2689_gather_scatter
    process(ptr_deref_2689_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2689_data_0;
      ov(31 downto 0) := iv;
      tmp28_2690 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2689_root_address_inst
    process(ptr_deref_2689_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2689_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2689_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2706_addr_0
    process(ptr_deref_2706_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2706_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2706_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2706_base_resize
    process(iNsTr_7_2703) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2703;
      ov := iv(0 downto 0);
      ptr_deref_2706_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2706_gather_scatter
    process(ptr_deref_2706_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2706_data_0;
      ov(15 downto 0) := iv;
      tmp36_2707 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2706_root_address_inst
    process(ptr_deref_2706_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2706_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2706_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2722_addr_0
    process(ptr_deref_2722_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2722_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2722_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2722_base_resize
    process(iNsTr_8_2719) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2719;
      ov := iv(6 downto 0);
      ptr_deref_2722_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2722_gather_scatter
    process(ptr_deref_2722_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2722_data_0;
      ov(31 downto 0) := iv;
      tmp39_2723 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2722_root_address_inst
    process(ptr_deref_2722_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2722_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2722_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2734_addr_0
    process(ptr_deref_2734_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2734_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2734_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2734_base_resize
    process(iNsTr_9_2731) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2731;
      ov := iv(6 downto 0);
      ptr_deref_2734_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2734_gather_scatter
    process(ptr_deref_2734_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2734_data_0;
      ov(31 downto 0) := iv;
      tmp48_2735 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2734_root_address_inst
    process(ptr_deref_2734_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2734_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2734_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2746_addr_0
    process(ptr_deref_2746_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2746_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2746_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2746_base_resize
    process(iNsTr_10_2743) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2743;
      ov := iv(6 downto 0);
      ptr_deref_2746_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2746_gather_scatter
    process(ptr_deref_2746_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2746_data_0;
      ov(31 downto 0) := iv;
      tmp51_2747 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2746_root_address_inst
    process(ptr_deref_2746_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2746_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2746_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2934_addr_0
    process(ptr_deref_2934_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2934_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2934_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2934_base_resize
    process(arrayidx_2931) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2931;
      ov := iv(13 downto 0);
      ptr_deref_2934_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2934_gather_scatter
    process(ptr_deref_2934_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2934_data_0;
      ov(63 downto 0) := iv;
      tmp61_2935 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2934_root_address_inst
    process(ptr_deref_2934_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2934_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2934_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2964_addr_0
    process(ptr_deref_2964_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2964_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2964_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2964_base_resize
    process(arrayidx66_2962) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx66_2962;
      ov := iv(13 downto 0);
      ptr_deref_2964_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2964_gather_scatter
    process(tmp61_2935) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp61_2935;
      ov(63 downto 0) := iv;
      ptr_deref_2964_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2964_root_address_inst
    process(ptr_deref_2964_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2964_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2964_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2983_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2982;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2983_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2983_branch_req_0,
          ack0 => if_stmt_2983_branch_ack_0,
          ack1 => if_stmt_2983_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3014_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp81_3013;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3014_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3014_branch_req_0,
          ack0 => if_stmt_3014_branch_ack_0,
          ack1 => if_stmt_3014_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3062_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp92_3061;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3062_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3062_branch_req_0,
          ack0 => if_stmt_3062_branch_ack_0,
          ack1 => if_stmt_3062_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2994_inst
    process(indvar_2877) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2877, type_cast_2993_wire_constant, tmp_var);
      indvarx_xnext_2995 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3002_inst
    process(input_dim1x_x1x_xph_2750) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2750, type_cast_3001_wire_constant, tmp_var);
      inc_3003 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3025_inst
    process(input_dim0x_x2x_xph_2756) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_2756, type_cast_3024_wire_constant, tmp_var);
      inc85_3026 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2781_inst
    process(mul_2777, conv16_2767) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_2777, conv16_2767, tmp_var);
      add_2782 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2796_inst
    process(mul27_2792, tmp28_2690) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul27_2792, tmp28_2690, tmp_var);
      add29_2797 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2811_inst
    process(mul38_2807, tmp39_2723) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul38_2807, tmp39_2723, tmp_var);
      add40_2812 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2828_inst
    process(sub44_2823) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub44_2823, type_cast_2827_wire_constant, tmp_var);
      sext_2829 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2849_inst
    process(sub32_2844) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub32_2844, type_cast_2848_wire_constant, tmp_var);
      sext106_2850 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2868_inst
    process(conv50_2838, mul54_2864) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv50_2838, mul54_2864, tmp_var);
      add55_2869 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2898_inst
    process(mul20_2787, conv13105_2894) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul20_2787, conv13105_2894, tmp_var);
      add21_2899 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2903_inst
    process(mul56_2874, conv13105_2894) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul56_2874, conv13105_2894, tmp_var);
      add57_2904 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2976_inst
    process(conv69_2971) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv69_2971, type_cast_2975_wire_constant, tmp_var);
      add70_2977 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2836_inst
    process(type_cast_2832_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2832_wire, type_cast_2835_wire_constant, tmp_var);
      ASHR_i32_i32_2836_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2857_inst
    process(type_cast_2853_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2853_wire, type_cast_2856_wire_constant, tmp_var);
      ASHR_i32_i32_2857_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2917_inst
    process(type_cast_2913_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2913_wire, type_cast_2916_wire_constant, tmp_var);
      ASHR_i32_i32_2917_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2948_inst
    process(type_cast_2944_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2944_wire, type_cast_2947_wire_constant, tmp_var);
      ASHR_i32_i32_2948_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3012_inst
    process(conv79_3008, tmp2_2642) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv79_3008, tmp2_2642, tmp_var);
      cmp81_3013 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3060_inst
    process(conv90_3056, tmp_2620) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv90_3056, tmp_2620, tmp_var);
      cmp92_3061 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2625_inst
    process(tmp_2620) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2620, type_cast_2624_wire_constant, tmp_var);
      div_2626 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2647_inst
    process(tmp2_2642) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp2_2642, type_cast_2646_wire_constant, tmp_var);
      div3_2648 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3031_inst
    process(tmp2_2642) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp2_2642, type_cast_3030_wire_constant, tmp_var);
      div87_3032 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2889_inst
    process(indvar_2877) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2877, type_cast_2888_wire_constant, tmp_var);
      input_dim2x_x1_2890 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2776_inst
    process(tmp2_2642, conv19_2772) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp2_2642, conv19_2772, tmp_var);
      mul_2777 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2786_inst
    process(add_2782, tmp14_2664) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_2782, tmp14_2664, tmp_var);
      mul20_2787 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2791_inst
    process(conv26_2678, conv19_2772) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv26_2678, conv19_2772, tmp_var);
      mul27_2792 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2806_inst
    process(conv37_2711, conv16_2767) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv37_2711, conv16_2767, tmp_var);
      mul38_2807 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2863_inst
    process(tmp51_2747, conv53_2859) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp51_2747, conv53_2859, tmp_var);
      mul54_2864 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2873_inst
    process(add55_2869, tmp48_2735) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add55_2869, tmp48_2735, tmp_var);
      mul56_2874 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2822_inst
    process(sub43_2817) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub43_2817, type_cast_2821_wire_constant, tmp_var);
      sub44_2823 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2843_inst
    process(sub_2802) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2802, type_cast_2842_wire_constant, tmp_var);
      sub32_2844 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2909_inst
    process(add21_2899) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add21_2899, type_cast_2908_wire_constant, tmp_var);
      sext108_2910 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2940_inst
    process(add57_2904) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add57_2904, type_cast_2939_wire_constant, tmp_var);
      sext109_2941 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2801_inst
    process(add29_2797, conv31_2697) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add29_2797, conv31_2697, tmp_var);
      sub_2802 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2816_inst
    process(add40_2812, conv31_2697) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add40_2812, conv31_2697, tmp_var);
      sub43_2817 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2981_inst
    process(add70_2977, tmp14_2664) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add70_2977, tmp14_2664, tmp_var);
      cmp_2982 <= tmp_var; --
    end process;
    -- shared split operator group (35) : array_obj_ref_2929_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2928_scaled;
      array_obj_ref_2929_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2929_index_offset_req_0;
      array_obj_ref_2929_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2929_index_offset_req_1;
      array_obj_ref_2929_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_2960_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom65_2959_scaled;
      array_obj_ref_2960_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2960_index_offset_req_0;
      array_obj_ref_2960_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2960_index_offset_req_1;
      array_obj_ref_2960_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- unary operator type_cast_2765_inst
    process(input_dim1x_x1x_xph_2750) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_2750, tmp_var);
      type_cast_2765_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2770_inst
    process(input_dim0x_x2x_xph_2756) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_2756, tmp_var);
      type_cast_2770_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2922_inst
    process(shr_2919) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2919, tmp_var);
      type_cast_2922_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2953_inst
    process(shr64_2950) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr64_2950, tmp_var);
      type_cast_2953_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2969_inst
    process(input_dim2x_x1_2890) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2890, tmp_var);
      type_cast_2969_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3006_inst
    process(inc_3003) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_3003, tmp_var);
      type_cast_3006_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3054_inst
    process(input_dim0x_x0_3045) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_3045, tmp_var);
      type_cast_3054_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_2692_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2692_load_0_req_0;
      LOAD_padding_2692_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2692_load_0_req_1;
      LOAD_padding_2692_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2692_word_address_0;
      LOAD_padding_2692_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2619_load_0 ptr_deref_2641_load_0 ptr_deref_2663_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2619_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2641_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2663_load_0_req_0;
      ptr_deref_2619_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2641_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2663_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2619_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2641_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2663_load_0_req_1;
      ptr_deref_2619_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2641_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2663_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2619_word_address_0 & ptr_deref_2641_word_address_0 & ptr_deref_2663_word_address_0;
      ptr_deref_2619_data_0 <= data_out(95 downto 64);
      ptr_deref_2641_data_0 <= data_out(63 downto 32);
      ptr_deref_2663_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2706_load_0 ptr_deref_2673_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2706_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2673_load_0_req_0;
      ptr_deref_2706_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2673_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2706_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2673_load_0_req_1;
      ptr_deref_2706_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2673_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2706_word_address_0 & ptr_deref_2673_word_address_0;
      ptr_deref_2706_data_0 <= data_out(31 downto 16);
      ptr_deref_2673_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2689_load_0 ptr_deref_2722_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2689_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2722_load_0_req_0;
      ptr_deref_2689_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2722_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2689_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2722_load_0_req_1;
      ptr_deref_2689_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2722_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2689_word_address_0 & ptr_deref_2722_word_address_0;
      ptr_deref_2689_data_0 <= data_out(63 downto 32);
      ptr_deref_2722_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2734_load_0 ptr_deref_2746_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2734_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2746_load_0_req_0;
      ptr_deref_2734_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2746_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2734_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2746_load_0_req_1;
      ptr_deref_2734_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2746_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2734_word_address_0 & ptr_deref_2746_word_address_0;
      ptr_deref_2734_data_0 <= data_out(63 downto 32);
      ptr_deref_2746_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2934_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2934_load_0_req_0;
      ptr_deref_2934_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2934_load_0_req_1;
      ptr_deref_2934_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2934_word_address_0;
      ptr_deref_2934_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2964_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2964_store_0_req_0;
      ptr_deref_2964_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2964_store_0_req_1;
      ptr_deref_2964_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2964_word_address_0;
      data_in <= ptr_deref_2964_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2606_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_start_2606_inst_req_0;
      RPIPE_Block3_start_2606_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_start_2606_inst_req_1;
      RPIPE_Block3_start_2606_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2607 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_3070_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_3070_inst_req_0;
      WPIPE_Block3_done_3070_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_3070_inst_req_1;
      WPIPE_Block3_done_3070_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2607;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_2864_start: Boolean;
  signal sendOutput_CP_2864_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_965_load_0_ack_0 : boolean;
  signal ptr_deref_965_load_0_req_0 : boolean;
  signal ptr_deref_965_load_0_req_1 : boolean;
  signal ptr_deref_965_load_0_ack_1 : boolean;
  signal ptr_deref_977_load_0_req_0 : boolean;
  signal ptr_deref_977_load_0_ack_0 : boolean;
  signal ptr_deref_977_load_0_req_1 : boolean;
  signal ptr_deref_977_load_0_ack_1 : boolean;
  signal ptr_deref_989_load_0_req_0 : boolean;
  signal ptr_deref_989_load_0_ack_0 : boolean;
  signal ptr_deref_989_load_0_req_1 : boolean;
  signal ptr_deref_989_load_0_ack_1 : boolean;
  signal type_cast_1003_inst_req_0 : boolean;
  signal type_cast_1003_inst_ack_0 : boolean;
  signal type_cast_1003_inst_req_1 : boolean;
  signal type_cast_1003_inst_ack_1 : boolean;
  signal if_stmt_1017_branch_req_0 : boolean;
  signal if_stmt_1017_branch_ack_1 : boolean;
  signal if_stmt_1017_branch_ack_0 : boolean;
  signal type_cast_1036_inst_req_0 : boolean;
  signal type_cast_1036_inst_ack_0 : boolean;
  signal type_cast_1036_inst_req_1 : boolean;
  signal type_cast_1036_inst_ack_1 : boolean;
  signal array_obj_ref_1071_index_offset_req_0 : boolean;
  signal array_obj_ref_1071_index_offset_ack_0 : boolean;
  signal array_obj_ref_1071_index_offset_req_1 : boolean;
  signal array_obj_ref_1071_index_offset_ack_1 : boolean;
  signal addr_of_1072_final_reg_req_0 : boolean;
  signal addr_of_1072_final_reg_ack_0 : boolean;
  signal addr_of_1072_final_reg_req_1 : boolean;
  signal addr_of_1072_final_reg_ack_1 : boolean;
  signal ptr_deref_1076_load_0_req_0 : boolean;
  signal ptr_deref_1076_load_0_ack_0 : boolean;
  signal ptr_deref_1076_load_0_req_1 : boolean;
  signal ptr_deref_1076_load_0_ack_1 : boolean;
  signal type_cast_1080_inst_req_0 : boolean;
  signal type_cast_1080_inst_ack_0 : boolean;
  signal type_cast_1080_inst_req_1 : boolean;
  signal type_cast_1080_inst_ack_1 : boolean;
  signal type_cast_1090_inst_req_0 : boolean;
  signal type_cast_1090_inst_ack_0 : boolean;
  signal type_cast_1090_inst_req_1 : boolean;
  signal type_cast_1090_inst_ack_1 : boolean;
  signal type_cast_1100_inst_req_0 : boolean;
  signal type_cast_1100_inst_ack_0 : boolean;
  signal type_cast_1100_inst_req_1 : boolean;
  signal type_cast_1100_inst_ack_1 : boolean;
  signal type_cast_1110_inst_req_0 : boolean;
  signal type_cast_1110_inst_ack_0 : boolean;
  signal type_cast_1110_inst_req_1 : boolean;
  signal type_cast_1110_inst_ack_1 : boolean;
  signal type_cast_1120_inst_req_0 : boolean;
  signal type_cast_1120_inst_ack_0 : boolean;
  signal type_cast_1120_inst_req_1 : boolean;
  signal type_cast_1120_inst_ack_1 : boolean;
  signal type_cast_1130_inst_req_0 : boolean;
  signal type_cast_1130_inst_ack_0 : boolean;
  signal type_cast_1130_inst_req_1 : boolean;
  signal type_cast_1130_inst_ack_1 : boolean;
  signal type_cast_1140_inst_req_0 : boolean;
  signal type_cast_1140_inst_ack_0 : boolean;
  signal type_cast_1140_inst_req_1 : boolean;
  signal type_cast_1140_inst_ack_1 : boolean;
  signal type_cast_1150_inst_req_0 : boolean;
  signal type_cast_1150_inst_ack_0 : boolean;
  signal type_cast_1150_inst_req_1 : boolean;
  signal type_cast_1150_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1152_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1152_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1152_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1152_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1155_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1155_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1155_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1155_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1158_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1158_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1158_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1158_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1161_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1161_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1161_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1161_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1164_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1164_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1164_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1164_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1167_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1167_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1167_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1167_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1170_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1170_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1170_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1170_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1173_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1173_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1173_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1173_inst_ack_1 : boolean;
  signal if_stmt_1187_branch_req_0 : boolean;
  signal if_stmt_1187_branch_ack_1 : boolean;
  signal if_stmt_1187_branch_ack_0 : boolean;
  signal phi_stmt_1059_req_0 : boolean;
  signal type_cast_1065_inst_req_0 : boolean;
  signal type_cast_1065_inst_ack_0 : boolean;
  signal type_cast_1065_inst_req_1 : boolean;
  signal type_cast_1065_inst_ack_1 : boolean;
  signal phi_stmt_1059_req_1 : boolean;
  signal phi_stmt_1059_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_2864_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_2864_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_2864_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_2864_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_2864: Block -- control-path 
    signal sendOutput_CP_2864_elements: BooleanArray(68 downto 0);
    -- 
  begin -- 
    sendOutput_CP_2864_elements(0) <= sendOutput_CP_2864_start;
    sendOutput_CP_2864_symbol <= sendOutput_CP_2864_elements(68);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	9 
    -- CP-element group 0:  members (86) 
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_update_start_
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_954/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/branch_block_stmt_954__entry__
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016__entry__
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_update_start_
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_update_start_
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/type_cast_1003_update_start_
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/type_cast_1003_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/type_cast_1003_Update/cr
      -- 
    rr_2927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(0), ack => ptr_deref_965_load_0_req_0); -- 
    cr_2938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(0), ack => ptr_deref_965_load_0_req_1); -- 
    rr_2977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(0), ack => ptr_deref_977_load_0_req_0); -- 
    cr_2988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(0), ack => ptr_deref_977_load_0_req_1); -- 
    rr_3027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(0), ack => ptr_deref_989_load_0_req_0); -- 
    cr_3038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(0), ack => ptr_deref_989_load_0_req_1); -- 
    cr_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(0), ack => type_cast_1003_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_sample_completed_
      -- 
    ra_2928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_965_load_0_ack_0, ack => sendOutput_CP_2864_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Update/ptr_deref_965_Merge/merge_ack
      -- CP-element group 2: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Update/ptr_deref_965_Merge/$exit
      -- CP-element group 2: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Update/ptr_deref_965_Merge/merge_req
      -- CP-element group 2: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_Update/ptr_deref_965_Merge/$entry
      -- CP-element group 2: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_965_update_completed_
      -- 
    ca_2939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_965_load_0_ack_1, ack => sendOutput_CP_2864_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Sample/word_access_start/word_0/ra
      -- 
    ra_2978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_977_load_0_ack_0, ack => sendOutput_CP_2864_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Update/ptr_deref_977_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Update/ptr_deref_977_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Update/ptr_deref_977_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_977_Update/ptr_deref_977_Merge/merge_ack
      -- 
    ca_2989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_977_load_0_ack_1, ack => sendOutput_CP_2864_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Sample/word_access_start/word_0/ra
      -- 
    ra_3028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_989_load_0_ack_0, ack => sendOutput_CP_2864_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Update/ptr_deref_989_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Update/ptr_deref_989_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Update/ptr_deref_989_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/ptr_deref_989_Update/ptr_deref_989_Merge/merge_ack
      -- 
    ca_3039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_989_load_0_ack_1, ack => sendOutput_CP_2864_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	6 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/type_cast_1003_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/type_cast_1003_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/type_cast_1003_Sample/rr
      -- 
    rr_3052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(7), ack => type_cast_1003_inst_req_0); -- 
    sendOutput_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "sendOutput_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_2864_elements(2) & sendOutput_CP_2864_elements(6) & sendOutput_CP_2864_elements(4);
      gj_sendOutput_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2864_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/type_cast_1003_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/type_cast_1003_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/type_cast_1003_Sample/ra
      -- 
    ra_3053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1003_inst_ack_0, ack => sendOutput_CP_2864_elements(8)); -- 
    -- CP-element group 9:  branch  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (13) 
      -- CP-element group 9: 	 branch_block_stmt_954/R_cmp77_1018_place
      -- CP-element group 9: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016__exit__
      -- CP-element group 9: 	 branch_block_stmt_954/if_stmt_1017__entry__
      -- CP-element group 9: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/$exit
      -- CP-element group 9: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/type_cast_1003_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/type_cast_1003_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_954/assign_stmt_962_to_assign_stmt_1016/type_cast_1003_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_954/if_stmt_1017_dead_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_954/if_stmt_1017_eval_test/$entry
      -- CP-element group 9: 	 branch_block_stmt_954/if_stmt_1017_eval_test/$exit
      -- CP-element group 9: 	 branch_block_stmt_954/if_stmt_1017_eval_test/branch_req
      -- CP-element group 9: 	 branch_block_stmt_954/if_stmt_1017_if_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_954/if_stmt_1017_else_link/$entry
      -- 
    ca_3058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1003_inst_ack_1, ack => sendOutput_CP_2864_elements(9)); -- 
    branch_req_3066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(9), ack => if_stmt_1017_branch_req_0); -- 
    -- CP-element group 10:  transition  place  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	68 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 branch_block_stmt_954/entry_forx_xend
      -- CP-element group 10: 	 branch_block_stmt_954/if_stmt_1017_if_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_954/if_stmt_1017_if_link/if_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_954/entry_forx_xend_PhiReq/$entry
      -- CP-element group 10: 	 branch_block_stmt_954/entry_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_3071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1017_branch_ack_1, ack => sendOutput_CP_2864_elements(10)); -- 
    -- CP-element group 11:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (18) 
      -- CP-element group 11: 	 branch_block_stmt_954/entry_bbx_xnph
      -- CP-element group 11: 	 branch_block_stmt_954/merge_stmt_1023__exit__
      -- CP-element group 11: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056__entry__
      -- CP-element group 11: 	 branch_block_stmt_954/if_stmt_1017_else_link/$exit
      -- CP-element group 11: 	 branch_block_stmt_954/if_stmt_1017_else_link/else_choice_transition
      -- CP-element group 11: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/$entry
      -- CP-element group 11: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/type_cast_1036_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/type_cast_1036_update_start_
      -- CP-element group 11: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/type_cast_1036_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/type_cast_1036_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/type_cast_1036_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/type_cast_1036_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_954/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 11: 	 branch_block_stmt_954/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 11: 	 branch_block_stmt_954/merge_stmt_1023_PhiReqMerge
      -- CP-element group 11: 	 branch_block_stmt_954/merge_stmt_1023_PhiAck/$entry
      -- CP-element group 11: 	 branch_block_stmt_954/merge_stmt_1023_PhiAck/$exit
      -- CP-element group 11: 	 branch_block_stmt_954/merge_stmt_1023_PhiAck/dummy
      -- 
    else_choice_transition_3075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1017_branch_ack_0, ack => sendOutput_CP_2864_elements(11)); -- 
    rr_3088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(11), ack => type_cast_1036_inst_req_0); -- 
    cr_3093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(11), ack => type_cast_1036_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/type_cast_1036_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/type_cast_1036_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/type_cast_1036_Sample/ra
      -- 
    ra_3089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1036_inst_ack_0, ack => sendOutput_CP_2864_elements(12)); -- 
    -- CP-element group 13:  transition  place  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	62 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056__exit__
      -- CP-element group 13: 	 branch_block_stmt_954/bbx_xnph_forx_xbody
      -- CP-element group 13: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/$exit
      -- CP-element group 13: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/type_cast_1036_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/type_cast_1036_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_954/assign_stmt_1028_to_assign_stmt_1056/type_cast_1036_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_954/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 13: 	 branch_block_stmt_954/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1059/$entry
      -- CP-element group 13: 	 branch_block_stmt_954/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/$entry
      -- 
    ca_3094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1036_inst_ack_1, ack => sendOutput_CP_2864_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	67 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	59 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_final_index_sum_regn_sample_complete
      -- CP-element group 14: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_final_index_sum_regn_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_final_index_sum_regn_Sample/ack
      -- 
    ack_3123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1071_index_offset_ack_0, ack => sendOutput_CP_2864_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	67 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (11) 
      -- CP-element group 15: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/addr_of_1072_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_offset_calculated
      -- CP-element group 15: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_final_index_sum_regn_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_final_index_sum_regn_Update/ack
      -- CP-element group 15: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/addr_of_1072_request/$entry
      -- CP-element group 15: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/addr_of_1072_request/req
      -- 
    ack_3128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1071_index_offset_ack_1, ack => sendOutput_CP_2864_elements(15)); -- 
    req_3137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(15), ack => addr_of_1072_final_reg_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/addr_of_1072_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/addr_of_1072_request/$exit
      -- CP-element group 16: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/addr_of_1072_request/ack
      -- 
    ack_3138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1072_final_reg_ack_0, ack => sendOutput_CP_2864_elements(16)); -- 
    -- CP-element group 17:  join  fork  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	67 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (24) 
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/addr_of_1072_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/addr_of_1072_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/addr_of_1072_complete/ack
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_base_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_word_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_root_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_base_address_resized
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_base_addr_resize/$entry
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_base_addr_resize/$exit
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_base_addr_resize/base_resize_req
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_base_addr_resize/base_resize_ack
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_base_plus_offset/$entry
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_base_plus_offset/$exit
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_base_plus_offset/sum_rename_req
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_base_plus_offset/sum_rename_ack
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_word_addrgen/$entry
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_word_addrgen/$exit
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_word_addrgen/root_register_req
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_word_addrgen/root_register_ack
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Sample/word_access_start/$entry
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Sample/word_access_start/word_0/$entry
      -- CP-element group 17: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Sample/word_access_start/word_0/rr
      -- 
    ack_3143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1072_final_reg_ack_1, ack => sendOutput_CP_2864_elements(17)); -- 
    rr_3176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(17), ack => ptr_deref_1076_load_0_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (5) 
      -- CP-element group 18: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Sample/word_access_start/$exit
      -- CP-element group 18: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Sample/word_access_start/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Sample/word_access_start/word_0/ra
      -- 
    ra_3177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1076_load_0_ack_0, ack => sendOutput_CP_2864_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	67 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	24 
    -- CP-element group 19: 	26 
    -- CP-element group 19: 	28 
    -- CP-element group 19: 	30 
    -- CP-element group 19: 	32 
    -- CP-element group 19: 	34 
    -- CP-element group 19:  members (33) 
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Update/word_access_complete/$exit
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Update/word_access_complete/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Update/word_access_complete/word_0/ca
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Update/ptr_deref_1076_Merge/$entry
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Update/ptr_deref_1076_Merge/$exit
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Update/ptr_deref_1076_Merge/merge_req
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Update/ptr_deref_1076_Merge/merge_ack
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1080_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1130_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1080_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1080_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1090_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1090_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1090_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1100_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1100_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1100_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1110_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1110_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1110_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1120_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1120_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1120_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1130_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1130_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1140_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1140_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1140_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1150_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1150_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1150_Sample/rr
      -- 
    ca_3188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1076_load_0_ack_1, ack => sendOutput_CP_2864_elements(19)); -- 
    rr_3201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(19), ack => type_cast_1080_inst_req_0); -- 
    rr_3215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(19), ack => type_cast_1090_inst_req_0); -- 
    rr_3229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(19), ack => type_cast_1100_inst_req_0); -- 
    rr_3243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(19), ack => type_cast_1110_inst_req_0); -- 
    rr_3257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(19), ack => type_cast_1120_inst_req_0); -- 
    rr_3271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(19), ack => type_cast_1130_inst_req_0); -- 
    rr_3285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(19), ack => type_cast_1140_inst_req_0); -- 
    rr_3299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(19), ack => type_cast_1150_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1080_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1080_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1080_Sample/ra
      -- 
    ra_3202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1080_inst_ack_0, ack => sendOutput_CP_2864_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	67 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	56 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1080_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1080_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1080_Update/ca
      -- 
    ca_3207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1080_inst_ack_1, ack => sendOutput_CP_2864_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1090_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1090_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1090_Sample/ra
      -- 
    ra_3216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1090_inst_ack_0, ack => sendOutput_CP_2864_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	67 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	53 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1090_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1090_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1090_Update/ca
      -- 
    ca_3221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1090_inst_ack_1, ack => sendOutput_CP_2864_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	19 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1100_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1100_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1100_Sample/ra
      -- 
    ra_3230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1100_inst_ack_0, ack => sendOutput_CP_2864_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	67 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	50 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1100_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1100_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1100_Update/ca
      -- 
    ca_3235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1100_inst_ack_1, ack => sendOutput_CP_2864_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	19 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1110_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1110_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1110_Sample/ra
      -- 
    ra_3244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_0, ack => sendOutput_CP_2864_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	67 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	47 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1110_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1110_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1110_Update/ca
      -- 
    ca_3249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_1, ack => sendOutput_CP_2864_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	19 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1120_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1120_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1120_Sample/ra
      -- 
    ra_3258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1120_inst_ack_0, ack => sendOutput_CP_2864_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	67 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	44 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1120_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1120_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1120_Update/ca
      -- 
    ca_3263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1120_inst_ack_1, ack => sendOutput_CP_2864_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	19 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1130_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1130_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1130_Sample/ra
      -- 
    ra_3272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1130_inst_ack_0, ack => sendOutput_CP_2864_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	67 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	41 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1130_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1130_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1130_Update/ca
      -- 
    ca_3277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1130_inst_ack_1, ack => sendOutput_CP_2864_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	19 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1140_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1140_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1140_Sample/ra
      -- 
    ra_3286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1140_inst_ack_0, ack => sendOutput_CP_2864_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	67 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	38 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1140_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1140_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1140_Update/ca
      -- 
    ca_3291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1140_inst_ack_1, ack => sendOutput_CP_2864_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	19 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1150_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1150_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1150_Sample/ra
      -- 
    ra_3300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1150_inst_ack_0, ack => sendOutput_CP_2864_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	67 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (6) 
      -- CP-element group 35: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1150_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1150_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1150_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1152_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1152_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1152_Sample/req
      -- 
    ca_3305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1150_inst_ack_1, ack => sendOutput_CP_2864_elements(35)); -- 
    req_3313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(35), ack => WPIPE_ConvTranspose_output_pipe_1152_inst_req_0); -- 
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1152_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1152_update_start_
      -- CP-element group 36: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1152_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1152_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1152_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1152_Update/req
      -- 
    ack_3314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1152_inst_ack_0, ack => sendOutput_CP_2864_elements(36)); -- 
    req_3318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(36), ack => WPIPE_ConvTranspose_output_pipe_1152_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1152_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1152_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1152_Update/ack
      -- 
    ack_3319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1152_inst_ack_1, ack => sendOutput_CP_2864_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	33 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1155_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1155_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1155_Sample/req
      -- 
    req_3327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(38), ack => WPIPE_ConvTranspose_output_pipe_1155_inst_req_0); -- 
    sendOutput_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2864_elements(33) & sendOutput_CP_2864_elements(37);
      gj_sendOutput_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2864_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1155_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1155_update_start_
      -- CP-element group 39: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1155_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1155_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1155_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1155_Update/req
      -- 
    ack_3328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1155_inst_ack_0, ack => sendOutput_CP_2864_elements(39)); -- 
    req_3332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(39), ack => WPIPE_ConvTranspose_output_pipe_1155_inst_req_1); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1155_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1155_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1155_Update/ack
      -- 
    ack_3333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1155_inst_ack_1, ack => sendOutput_CP_2864_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	31 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1158_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1158_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1158_Sample/req
      -- 
    req_3341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(41), ack => WPIPE_ConvTranspose_output_pipe_1158_inst_req_0); -- 
    sendOutput_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2864_elements(31) & sendOutput_CP_2864_elements(40);
      gj_sendOutput_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2864_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1158_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1158_update_start_
      -- CP-element group 42: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1158_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1158_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1158_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1158_Update/req
      -- 
    ack_3342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1158_inst_ack_0, ack => sendOutput_CP_2864_elements(42)); -- 
    req_3346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(42), ack => WPIPE_ConvTranspose_output_pipe_1158_inst_req_1); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1158_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1158_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1158_Update/ack
      -- 
    ack_3347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1158_inst_ack_1, ack => sendOutput_CP_2864_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	29 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1161_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1161_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1161_Sample/req
      -- 
    req_3355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(44), ack => WPIPE_ConvTranspose_output_pipe_1161_inst_req_0); -- 
    sendOutput_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2864_elements(29) & sendOutput_CP_2864_elements(43);
      gj_sendOutput_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2864_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1161_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1161_update_start_
      -- CP-element group 45: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1161_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1161_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1161_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1161_Update/req
      -- 
    ack_3356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1161_inst_ack_0, ack => sendOutput_CP_2864_elements(45)); -- 
    req_3360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(45), ack => WPIPE_ConvTranspose_output_pipe_1161_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1161_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1161_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1161_Update/ack
      -- 
    ack_3361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1161_inst_ack_1, ack => sendOutput_CP_2864_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	27 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1164_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1164_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1164_Sample/req
      -- 
    req_3369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(47), ack => WPIPE_ConvTranspose_output_pipe_1164_inst_req_0); -- 
    sendOutput_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2864_elements(27) & sendOutput_CP_2864_elements(46);
      gj_sendOutput_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2864_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1164_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1164_update_start_
      -- CP-element group 48: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1164_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1164_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1164_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1164_Update/req
      -- 
    ack_3370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1164_inst_ack_0, ack => sendOutput_CP_2864_elements(48)); -- 
    req_3374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(48), ack => WPIPE_ConvTranspose_output_pipe_1164_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1164_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1164_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1164_Update/ack
      -- 
    ack_3375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1164_inst_ack_1, ack => sendOutput_CP_2864_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	25 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1167_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1167_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1167_Sample/req
      -- 
    req_3383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(50), ack => WPIPE_ConvTranspose_output_pipe_1167_inst_req_0); -- 
    sendOutput_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2864_elements(25) & sendOutput_CP_2864_elements(49);
      gj_sendOutput_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2864_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1167_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1167_update_start_
      -- CP-element group 51: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1167_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1167_Sample/ack
      -- CP-element group 51: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1167_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1167_Update/req
      -- 
    ack_3384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1167_inst_ack_0, ack => sendOutput_CP_2864_elements(51)); -- 
    req_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(51), ack => WPIPE_ConvTranspose_output_pipe_1167_inst_req_1); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1167_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1167_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1167_Update/ack
      -- 
    ack_3389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1167_inst_ack_1, ack => sendOutput_CP_2864_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	23 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1170_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1170_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1170_Sample/req
      -- 
    req_3397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(53), ack => WPIPE_ConvTranspose_output_pipe_1170_inst_req_0); -- 
    sendOutput_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2864_elements(23) & sendOutput_CP_2864_elements(52);
      gj_sendOutput_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2864_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1170_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1170_update_start_
      -- CP-element group 54: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1170_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1170_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1170_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1170_Update/req
      -- 
    ack_3398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1170_inst_ack_0, ack => sendOutput_CP_2864_elements(54)); -- 
    req_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(54), ack => WPIPE_ConvTranspose_output_pipe_1170_inst_req_1); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1170_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1170_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1170_Update/ack
      -- 
    ack_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1170_inst_ack_1, ack => sendOutput_CP_2864_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	21 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1173_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1173_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1173_Sample/req
      -- 
    req_3411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(56), ack => WPIPE_ConvTranspose_output_pipe_1173_inst_req_0); -- 
    sendOutput_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2864_elements(21) & sendOutput_CP_2864_elements(55);
      gj_sendOutput_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2864_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1173_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1173_update_start_
      -- CP-element group 57: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1173_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1173_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1173_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1173_Update/req
      -- 
    ack_3412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1173_inst_ack_0, ack => sendOutput_CP_2864_elements(57)); -- 
    req_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(57), ack => WPIPE_ConvTranspose_output_pipe_1173_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1173_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1173_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/WPIPE_ConvTranspose_output_pipe_1173_Update/ack
      -- 
    ack_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1173_inst_ack_1, ack => sendOutput_CP_2864_elements(58)); -- 
    -- CP-element group 59:  branch  join  transition  place  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	14 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (10) 
      -- CP-element group 59: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186__exit__
      -- CP-element group 59: 	 branch_block_stmt_954/if_stmt_1187__entry__
      -- CP-element group 59: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/$exit
      -- CP-element group 59: 	 branch_block_stmt_954/if_stmt_1187_dead_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_954/if_stmt_1187_eval_test/$entry
      -- CP-element group 59: 	 branch_block_stmt_954/if_stmt_1187_eval_test/$exit
      -- CP-element group 59: 	 branch_block_stmt_954/if_stmt_1187_eval_test/branch_req
      -- CP-element group 59: 	 branch_block_stmt_954/R_exitcond9_1188_place
      -- CP-element group 59: 	 branch_block_stmt_954/if_stmt_1187_if_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_954/if_stmt_1187_else_link/$entry
      -- 
    branch_req_3425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(59), ack => if_stmt_1187_branch_req_0); -- 
    sendOutput_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2864_elements(14) & sendOutput_CP_2864_elements(58);
      gj_sendOutput_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2864_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  merge  transition  place  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	68 
    -- CP-element group 60:  members (13) 
      -- CP-element group 60: 	 branch_block_stmt_954/merge_stmt_1193__exit__
      -- CP-element group 60: 	 branch_block_stmt_954/forx_xendx_xloopexit_forx_xend
      -- CP-element group 60: 	 branch_block_stmt_954/if_stmt_1187_if_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_954/if_stmt_1187_if_link/if_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_954/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 60: 	 branch_block_stmt_954/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_954/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_954/merge_stmt_1193_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_954/merge_stmt_1193_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_954/merge_stmt_1193_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_954/merge_stmt_1193_PhiAck/dummy
      -- CP-element group 60: 	 branch_block_stmt_954/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_954/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_3430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1187_branch_ack_1, ack => sendOutput_CP_2864_elements(60)); -- 
    -- CP-element group 61:  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: 	64 
    -- CP-element group 61:  members (12) 
      -- CP-element group 61: 	 branch_block_stmt_954/if_stmt_1187_else_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_954/if_stmt_1187_else_link/else_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_954/forx_xbody_forx_xbody
      -- CP-element group 61: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/$entry
      -- CP-element group 61: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/$entry
      -- CP-element group 61: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1187_branch_ack_0, ack => sendOutput_CP_2864_elements(61)); -- 
    rr_3478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(61), ack => type_cast_1065_inst_req_0); -- 
    cr_3483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(61), ack => type_cast_1065_inst_req_1); -- 
    -- CP-element group 62:  transition  output  delay-element  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	13 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	66 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_954/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_954/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1059/$exit
      -- CP-element group 62: 	 branch_block_stmt_954/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/$exit
      -- CP-element group 62: 	 branch_block_stmt_954/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1063_konst_delay_trans
      -- CP-element group 62: 	 branch_block_stmt_954/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_req
      -- 
    phi_stmt_1059_req_3459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1059_req_3459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(62), ack => phi_stmt_1059_req_0); -- 
    -- Element group sendOutput_CP_2864_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => sendOutput_CP_2864_elements(13), ack => sendOutput_CP_2864_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Sample/ra
      -- 
    ra_3479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1065_inst_ack_0, ack => sendOutput_CP_2864_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	61 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Update/ca
      -- 
    ca_3484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1065_inst_ack_1, ack => sendOutput_CP_2864_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/$exit
      -- CP-element group 65: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/$exit
      -- CP-element group 65: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/$exit
      -- CP-element group 65: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/$exit
      -- CP-element group 65: 	 branch_block_stmt_954/forx_xbody_forx_xbody_PhiReq/phi_stmt_1059/phi_stmt_1059_req
      -- 
    phi_stmt_1059_req_3485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1059_req_3485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(65), ack => phi_stmt_1059_req_1); -- 
    sendOutput_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2864_elements(63) & sendOutput_CP_2864_elements(64);
      gj_sendOutput_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2864_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  merge  transition  place  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	62 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_954/merge_stmt_1058_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_954/merge_stmt_1058_PhiAck/$entry
      -- 
    sendOutput_CP_2864_elements(66) <= OrReduce(sendOutput_CP_2864_elements(62) & sendOutput_CP_2864_elements(65));
    -- CP-element group 67:  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	14 
    -- CP-element group 67: 	15 
    -- CP-element group 67: 	17 
    -- CP-element group 67: 	19 
    -- CP-element group 67: 	21 
    -- CP-element group 67: 	23 
    -- CP-element group 67: 	25 
    -- CP-element group 67: 	27 
    -- CP-element group 67: 	29 
    -- CP-element group 67: 	31 
    -- CP-element group 67: 	33 
    -- CP-element group 67: 	35 
    -- CP-element group 67:  members (53) 
      -- CP-element group 67: 	 branch_block_stmt_954/merge_stmt_1058__exit__
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186__entry__
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/addr_of_1072_update_start_
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_index_resized_1
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_index_scaled_1
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_index_computed_1
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_index_resize_1/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_index_resize_1/$exit
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_index_resize_1/index_resize_req
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_index_resize_1/index_resize_ack
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_index_scale_1/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_index_scale_1/$exit
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_index_scale_1/scale_rename_req
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_index_scale_1/scale_rename_ack
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_final_index_sum_regn_update_start
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_final_index_sum_regn_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_final_index_sum_regn_Sample/req
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_final_index_sum_regn_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/array_obj_ref_1071_final_index_sum_regn_Update/req
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/addr_of_1072_complete/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/addr_of_1072_complete/req
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_update_start_
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Update/word_access_complete/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Update/word_access_complete/word_0/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/ptr_deref_1076_Update/word_access_complete/word_0/cr
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1080_update_start_
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1080_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1080_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1090_update_start_
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1090_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1090_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1100_update_start_
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1100_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1100_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1110_update_start_
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1110_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1110_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1120_update_start_
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1120_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1120_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1130_update_start_
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1130_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1130_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1140_update_start_
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1140_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1140_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1150_update_start_
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1150_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_954/assign_stmt_1073_to_assign_stmt_1186/type_cast_1150_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_954/merge_stmt_1058_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_954/merge_stmt_1058_PhiAck/phi_stmt_1059_ack
      -- 
    phi_stmt_1059_ack_3490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1059_ack_0, ack => sendOutput_CP_2864_elements(67)); -- 
    req_3122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(67), ack => array_obj_ref_1071_index_offset_req_0); -- 
    req_3127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(67), ack => array_obj_ref_1071_index_offset_req_1); -- 
    req_3142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(67), ack => addr_of_1072_final_reg_req_1); -- 
    cr_3187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(67), ack => ptr_deref_1076_load_0_req_1); -- 
    cr_3206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(67), ack => type_cast_1080_inst_req_1); -- 
    cr_3220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(67), ack => type_cast_1090_inst_req_1); -- 
    cr_3234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(67), ack => type_cast_1100_inst_req_1); -- 
    cr_3248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(67), ack => type_cast_1110_inst_req_1); -- 
    cr_3262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(67), ack => type_cast_1120_inst_req_1); -- 
    cr_3276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(67), ack => type_cast_1130_inst_req_1); -- 
    cr_3290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(67), ack => type_cast_1140_inst_req_1); -- 
    cr_3304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2864_elements(67), ack => type_cast_1150_inst_req_1); -- 
    -- CP-element group 68:  merge  transition  place  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	10 
    -- CP-element group 68: 	60 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 $exit
      -- CP-element group 68: 	 branch_block_stmt_954/$exit
      -- CP-element group 68: 	 branch_block_stmt_954/branch_block_stmt_954__exit__
      -- CP-element group 68: 	 branch_block_stmt_954/merge_stmt_1195__exit__
      -- CP-element group 68: 	 branch_block_stmt_954/return__
      -- CP-element group 68: 	 branch_block_stmt_954/merge_stmt_1197__exit__
      -- CP-element group 68: 	 branch_block_stmt_954/merge_stmt_1195_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_954/merge_stmt_1195_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_954/merge_stmt_1195_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_954/merge_stmt_1195_PhiAck/dummy
      -- CP-element group 68: 	 branch_block_stmt_954/return___PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_954/return___PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_954/merge_stmt_1197_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_954/merge_stmt_1197_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_954/merge_stmt_1197_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_954/merge_stmt_1197_PhiAck/dummy
      -- 
    sendOutput_CP_2864_elements(68) <= OrReduce(sendOutput_CP_2864_elements(10) & sendOutput_CP_2864_elements(60));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_1070_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1070_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_1071_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1071_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1071_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1071_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1071_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1071_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_1073 : std_logic_vector(31 downto 0);
    signal cmp77_1016 : std_logic_vector(0 downto 0);
    signal conv14_1081 : std_logic_vector(7 downto 0);
    signal conv20_1091 : std_logic_vector(7 downto 0);
    signal conv26_1101 : std_logic_vector(7 downto 0);
    signal conv32_1111 : std_logic_vector(7 downto 0);
    signal conv38_1121 : std_logic_vector(7 downto 0);
    signal conv44_1131 : std_logic_vector(7 downto 0);
    signal conv50_1141 : std_logic_vector(7 downto 0);
    signal conv56_1151 : std_logic_vector(7 downto 0);
    signal conv_1004 : std_logic_vector(63 downto 0);
    signal exitcond9_1186 : std_logic_vector(0 downto 0);
    signal iNsTr_0_962 : std_logic_vector(31 downto 0);
    signal iNsTr_1_974 : std_logic_vector(31 downto 0);
    signal iNsTr_2_986 : std_logic_vector(31 downto 0);
    signal indvar_1059 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1181 : std_logic_vector(63 downto 0);
    signal mul3_1000 : std_logic_vector(31 downto 0);
    signal mul_995 : std_logic_vector(31 downto 0);
    signal ptr_deref_1076_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1076_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1076_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1076_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1076_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_965_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_965_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_965_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_965_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_965_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_977_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_977_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_977_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_977_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_977_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_989_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_989_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_989_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_989_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_989_word_offset_0 : std_logic_vector(6 downto 0);
    signal shr17_1087 : std_logic_vector(63 downto 0);
    signal shr23_1097 : std_logic_vector(63 downto 0);
    signal shr29_1107 : std_logic_vector(63 downto 0);
    signal shr35_1117 : std_logic_vector(63 downto 0);
    signal shr41_1127 : std_logic_vector(63 downto 0);
    signal shr47_1137 : std_logic_vector(63 downto 0);
    signal shr53_1147 : std_logic_vector(63 downto 0);
    signal shr76x_xmask_1010 : std_logic_vector(63 downto 0);
    signal tmp11_1077 : std_logic_vector(63 downto 0);
    signal tmp1_978 : std_logic_vector(31 downto 0);
    signal tmp2_990 : std_logic_vector(31 downto 0);
    signal tmp3_1028 : std_logic_vector(31 downto 0);
    signal tmp4_1033 : std_logic_vector(31 downto 0);
    signal tmp5_1037 : std_logic_vector(63 downto 0);
    signal tmp6_1043 : std_logic_vector(63 downto 0);
    signal tmp7_1049 : std_logic_vector(0 downto 0);
    signal tmp_966 : std_logic_vector(31 downto 0);
    signal type_cast_1008_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1014_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1041_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1047_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1054_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1063_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1065_wire : std_logic_vector(63 downto 0);
    signal type_cast_1085_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1095_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1105_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1115_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1125_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1135_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1145_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1179_wire_constant : std_logic_vector(63 downto 0);
    signal umax8_1056 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1071_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1071_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1071_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1071_resized_base_address <= "00000000000000";
    iNsTr_0_962 <= "00000000000000000000000000000010";
    iNsTr_1_974 <= "00000000000000000000000000000011";
    iNsTr_2_986 <= "00000000000000000000000000000100";
    ptr_deref_1076_word_offset_0 <= "00000000000000";
    ptr_deref_965_word_offset_0 <= "0000000";
    ptr_deref_977_word_offset_0 <= "0000000";
    ptr_deref_989_word_offset_0 <= "0000000";
    type_cast_1008_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_1014_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1041_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1047_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1054_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1063_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1085_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1095_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1105_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1115_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1125_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1135_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1145_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1179_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1059: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1063_wire_constant & type_cast_1065_wire;
      req <= phi_stmt_1059_req_0 & phi_stmt_1059_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1059",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1059_ack_0,
          idata => idata,
          odata => indvar_1059,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1059
    -- flow-through select operator MUX_1055_inst
    umax8_1056 <= tmp6_1043 when (tmp7_1049(0) /=  '0') else type_cast_1054_wire_constant;
    addr_of_1072_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1072_final_reg_req_0;
      addr_of_1072_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1072_final_reg_req_1;
      addr_of_1072_final_reg_ack_1<= rack(0);
      addr_of_1072_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1072_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1071_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1073,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1003_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1003_inst_req_0;
      type_cast_1003_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1003_inst_req_1;
      type_cast_1003_inst_ack_1<= rack(0);
      type_cast_1003_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1003_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul3_1000,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1004,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1036_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1036_inst_req_0;
      type_cast_1036_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1036_inst_req_1;
      type_cast_1036_inst_ack_1<= rack(0);
      type_cast_1036_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1036_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_1033,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp5_1037,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1065_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1065_inst_req_0;
      type_cast_1065_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1065_inst_req_1;
      type_cast_1065_inst_ack_1<= rack(0);
      type_cast_1065_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1065_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1181,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1065_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1080_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1080_inst_req_0;
      type_cast_1080_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1080_inst_req_1;
      type_cast_1080_inst_ack_1<= rack(0);
      type_cast_1080_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1080_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp11_1077,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv14_1081,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1090_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1090_inst_req_0;
      type_cast_1090_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1090_inst_req_1;
      type_cast_1090_inst_ack_1<= rack(0);
      type_cast_1090_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1090_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr17_1087,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_1091,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1100_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1100_inst_req_0;
      type_cast_1100_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1100_inst_req_1;
      type_cast_1100_inst_ack_1<= rack(0);
      type_cast_1100_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1100_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr23_1097,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_1101,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1110_inst_req_0;
      type_cast_1110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1110_inst_req_1;
      type_cast_1110_inst_ack_1<= rack(0);
      type_cast_1110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr29_1107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_1111,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1120_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1120_inst_req_0;
      type_cast_1120_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1120_inst_req_1;
      type_cast_1120_inst_ack_1<= rack(0);
      type_cast_1120_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1120_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr35_1117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_1121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1130_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1130_inst_req_0;
      type_cast_1130_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1130_inst_req_1;
      type_cast_1130_inst_ack_1<= rack(0);
      type_cast_1130_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1130_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr41_1127,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_1131,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1140_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1140_inst_req_0;
      type_cast_1140_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1140_inst_req_1;
      type_cast_1140_inst_ack_1<= rack(0);
      type_cast_1140_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1140_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr47_1137,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_1141,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1150_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1150_inst_req_0;
      type_cast_1150_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1150_inst_req_1;
      type_cast_1150_inst_ack_1<= rack(0);
      type_cast_1150_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1150_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr53_1147,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_1151,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1071_index_1_rename
    process(R_indvar_1070_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1070_resized;
      ov(13 downto 0) := iv;
      R_indvar_1070_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1071_index_1_resize
    process(indvar_1059) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1059;
      ov := iv(13 downto 0);
      R_indvar_1070_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1071_root_address_inst
    process(array_obj_ref_1071_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1071_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1071_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1076_addr_0
    process(ptr_deref_1076_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1076_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1076_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1076_base_resize
    process(arrayidx_1073) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1073;
      ov := iv(13 downto 0);
      ptr_deref_1076_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1076_gather_scatter
    process(ptr_deref_1076_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1076_data_0;
      ov(63 downto 0) := iv;
      tmp11_1077 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1076_root_address_inst
    process(ptr_deref_1076_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1076_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1076_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_965_addr_0
    process(ptr_deref_965_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_965_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_965_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_965_base_resize
    process(iNsTr_0_962) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_962;
      ov := iv(6 downto 0);
      ptr_deref_965_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_965_gather_scatter
    process(ptr_deref_965_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_965_data_0;
      ov(31 downto 0) := iv;
      tmp_966 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_965_root_address_inst
    process(ptr_deref_965_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_965_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_965_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_977_addr_0
    process(ptr_deref_977_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_977_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_977_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_977_base_resize
    process(iNsTr_1_974) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_974;
      ov := iv(6 downto 0);
      ptr_deref_977_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_977_gather_scatter
    process(ptr_deref_977_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_977_data_0;
      ov(31 downto 0) := iv;
      tmp1_978 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_977_root_address_inst
    process(ptr_deref_977_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_977_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_977_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_989_addr_0
    process(ptr_deref_989_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_989_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_989_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_989_base_resize
    process(iNsTr_2_986) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_986;
      ov := iv(6 downto 0);
      ptr_deref_989_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_989_gather_scatter
    process(ptr_deref_989_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_989_data_0;
      ov(31 downto 0) := iv;
      tmp2_990 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_989_root_address_inst
    process(ptr_deref_989_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_989_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_989_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_1017_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_1016;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1017_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1017_branch_req_0,
          ack0 => if_stmt_1017_branch_ack_0,
          ack1 => if_stmt_1017_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1187_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond9_1186;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1187_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1187_branch_req_0,
          ack0 => if_stmt_1187_branch_ack_0,
          ack1 => if_stmt_1187_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_1180_inst
    process(indvar_1059) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1059, type_cast_1179_wire_constant, tmp_var);
      indvarx_xnext_1181 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1009_inst
    process(conv_1004) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv_1004, type_cast_1008_wire_constant, tmp_var);
      shr76x_xmask_1010 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1015_inst
    process(shr76x_xmask_1010) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr76x_xmask_1010, type_cast_1014_wire_constant, tmp_var);
      cmp77_1016 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1185_inst
    process(indvarx_xnext_1181, umax8_1056) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1181, umax8_1056, tmp_var);
      exitcond9_1186 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1042_inst
    process(tmp5_1037) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_1037, type_cast_1041_wire_constant, tmp_var);
      tmp6_1043 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1086_inst
    process(tmp11_1077) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_1077, type_cast_1085_wire_constant, tmp_var);
      shr17_1087 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1096_inst
    process(tmp11_1077) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_1077, type_cast_1095_wire_constant, tmp_var);
      shr23_1097 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1106_inst
    process(tmp11_1077) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_1077, type_cast_1105_wire_constant, tmp_var);
      shr29_1107 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1116_inst
    process(tmp11_1077) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_1077, type_cast_1115_wire_constant, tmp_var);
      shr35_1117 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1126_inst
    process(tmp11_1077) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_1077, type_cast_1125_wire_constant, tmp_var);
      shr41_1127 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1136_inst
    process(tmp11_1077) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_1077, type_cast_1135_wire_constant, tmp_var);
      shr47_1137 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1146_inst
    process(tmp11_1077) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_1077, type_cast_1145_wire_constant, tmp_var);
      shr53_1147 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1027_inst
    process(tmp1_978, tmp_966) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_978, tmp_966, tmp_var);
      tmp3_1028 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1032_inst
    process(tmp3_1028, tmp2_990) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp3_1028, tmp2_990, tmp_var);
      tmp4_1033 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_994_inst
    process(tmp1_978, tmp_966) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_978, tmp_966, tmp_var);
      mul_995 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_999_inst
    process(mul_995, tmp2_990) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_995, tmp2_990, tmp_var);
      mul3_1000 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1048_inst
    process(tmp6_1043) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp6_1043, type_cast_1047_wire_constant, tmp_var);
      tmp7_1049 <= tmp_var; --
    end process;
    -- shared split operator group (17) : array_obj_ref_1071_index_offset 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1070_scaled;
      array_obj_ref_1071_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1071_index_offset_req_0;
      array_obj_ref_1071_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1071_index_offset_req_1;
      array_obj_ref_1071_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_17_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared load operator group (0) : ptr_deref_1076_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1076_load_0_req_0;
      ptr_deref_1076_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1076_load_0_req_1;
      ptr_deref_1076_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1076_word_address_0;
      ptr_deref_1076_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(13 downto 0),
          mtag => memory_space_5_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(63 downto 0),
          mtag => memory_space_5_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_989_load_0 ptr_deref_977_load_0 ptr_deref_965_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_989_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_977_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_965_load_0_req_0;
      ptr_deref_989_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_977_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_965_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_989_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_977_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_965_load_0_req_1;
      ptr_deref_989_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_977_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_965_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_989_word_address_0 & ptr_deref_977_word_address_0 & ptr_deref_965_word_address_0;
      ptr_deref_989_data_0 <= data_out(95 downto 64);
      ptr_deref_977_data_0 <= data_out(63 downto 32);
      ptr_deref_965_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared outport operator group (0) : WPIPE_ConvTranspose_output_pipe_1173_inst WPIPE_ConvTranspose_output_pipe_1158_inst WPIPE_ConvTranspose_output_pipe_1152_inst WPIPE_ConvTranspose_output_pipe_1161_inst WPIPE_ConvTranspose_output_pipe_1164_inst WPIPE_ConvTranspose_output_pipe_1170_inst WPIPE_ConvTranspose_output_pipe_1167_inst WPIPE_ConvTranspose_output_pipe_1155_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1173_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1158_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1152_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1161_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1164_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1170_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1167_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1155_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1173_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1158_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1152_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1161_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1164_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1170_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1167_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1155_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1173_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1158_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1152_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1161_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1164_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1170_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1167_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1155_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1173_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1158_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1152_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1161_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1164_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1170_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1167_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1155_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv14_1081 & conv44_1131 & conv56_1151 & conv38_1121 & conv32_1111 & conv20_1091 & conv26_1101 & conv50_1141;
      ConvTranspose_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal ret_val_x_x_update_enable: Boolean;
  signal testConfigure_CP_0_start: Boolean;
  signal testConfigure_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal if_stmt_500_branch_req_0 : boolean;
  signal ptr_deref_405_load_0_req_1 : boolean;
  signal type_cast_83_inst_req_0 : boolean;
  signal if_stmt_936_branch_ack_1 : boolean;
  signal if_stmt_500_branch_ack_0 : boolean;
  signal if_stmt_500_branch_ack_1 : boolean;
  signal type_cast_486_inst_ack_0 : boolean;
  signal type_cast_947_inst_ack_0 : boolean;
  signal ptr_deref_368_store_0_req_1 : boolean;
  signal ptr_deref_368_store_0_ack_0 : boolean;
  signal ptr_deref_368_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 : boolean;
  signal type_cast_947_inst_ack_1 : boolean;
  signal type_cast_38_inst_req_0 : boolean;
  signal type_cast_38_inst_ack_0 : boolean;
  signal type_cast_38_inst_req_1 : boolean;
  signal type_cast_38_inst_ack_1 : boolean;
  signal type_cast_267_inst_req_1 : boolean;
  signal ptr_deref_405_load_0_req_0 : boolean;
  signal ptr_deref_455_load_0_ack_1 : boolean;
  signal ptr_deref_122_load_0_req_0 : boolean;
  signal ptr_deref_122_load_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_874_inst_ack_0 : boolean;
  signal ptr_deref_47_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_910_inst_ack_0 : boolean;
  signal ptr_deref_47_store_0_ack_0 : boolean;
  signal phi_stmt_73_req_1 : boolean;
  signal ptr_deref_47_store_0_req_1 : boolean;
  signal ptr_deref_47_store_0_ack_1 : boolean;
  signal type_cast_357_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_ack_0 : boolean;
  signal type_cast_896_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_ack_1 : boolean;
  signal type_cast_153_inst_req_0 : boolean;
  signal type_cast_947_inst_req_0 : boolean;
  signal type_cast_62_inst_req_0 : boolean;
  signal type_cast_62_inst_ack_0 : boolean;
  signal type_cast_62_inst_req_1 : boolean;
  signal type_cast_62_inst_ack_1 : boolean;
  signal ptr_deref_443_load_0_ack_1 : boolean;
  signal if_stmt_64_branch_req_0 : boolean;
  signal if_stmt_64_branch_ack_1 : boolean;
  signal type_cast_83_inst_req_1 : boolean;
  signal if_stmt_64_branch_ack_0 : boolean;
  signal type_cast_486_inst_req_0 : boolean;
  signal ptr_deref_443_load_0_req_1 : boolean;
  signal type_cast_95_inst_req_0 : boolean;
  signal type_cast_914_inst_req_0 : boolean;
  signal type_cast_95_inst_ack_0 : boolean;
  signal type_cast_95_inst_req_1 : boolean;
  signal type_cast_357_inst_req_1 : boolean;
  signal type_cast_95_inst_ack_1 : boolean;
  signal if_stmt_936_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_856_inst_req_0 : boolean;
  signal ptr_deref_431_load_0_ack_1 : boolean;
  signal ptr_deref_431_load_0_req_1 : boolean;
  signal array_obj_ref_101_index_offset_req_0 : boolean;
  signal array_obj_ref_101_index_offset_ack_0 : boolean;
  signal array_obj_ref_101_index_offset_req_1 : boolean;
  signal array_obj_ref_101_index_offset_ack_1 : boolean;
  signal ptr_deref_467_load_0_ack_1 : boolean;
  signal type_cast_153_inst_ack_0 : boolean;
  signal addr_of_102_final_reg_req_0 : boolean;
  signal addr_of_102_final_reg_ack_0 : boolean;
  signal addr_of_102_final_reg_req_1 : boolean;
  signal addr_of_102_final_reg_ack_1 : boolean;
  signal type_cast_914_inst_ack_0 : boolean;
  signal type_cast_419_inst_ack_1 : boolean;
  signal ptr_deref_405_load_0_ack_0 : boolean;
  signal type_cast_419_inst_req_1 : boolean;
  signal ptr_deref_105_store_0_req_0 : boolean;
  signal ptr_deref_105_store_0_ack_0 : boolean;
  signal ptr_deref_105_store_0_req_1 : boolean;
  signal ptr_deref_105_store_0_ack_1 : boolean;
  signal ptr_deref_431_load_0_ack_0 : boolean;
  signal ptr_deref_431_load_0_req_0 : boolean;
  signal type_cast_153_inst_req_1 : boolean;
  signal phi_stmt_264_req_0 : boolean;
  signal ptr_deref_381_load_0_ack_0 : boolean;
  signal ptr_deref_277_store_0_req_0 : boolean;
  signal ptr_deref_122_load_0_req_1 : boolean;
  signal ptr_deref_122_load_0_ack_1 : boolean;
  signal ptr_deref_455_load_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_130_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_130_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_130_inst_req_1 : boolean;
  signal type_cast_419_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_130_inst_ack_1 : boolean;
  signal type_cast_134_inst_req_0 : boolean;
  signal type_cast_134_inst_ack_0 : boolean;
  signal type_cast_134_inst_req_1 : boolean;
  signal type_cast_419_inst_req_0 : boolean;
  signal type_cast_134_inst_ack_1 : boolean;
  signal ptr_deref_467_load_0_req_1 : boolean;
  signal type_cast_83_inst_ack_1 : boolean;
  signal if_stmt_136_branch_req_0 : boolean;
  signal type_cast_357_inst_ack_0 : boolean;
  signal ptr_deref_443_load_0_ack_0 : boolean;
  signal if_stmt_136_branch_ack_1 : boolean;
  signal if_stmt_136_branch_ack_0 : boolean;
  signal type_cast_153_inst_ack_1 : boolean;
  signal ptr_deref_443_load_0_req_0 : boolean;
  signal ptr_deref_164_store_0_req_0 : boolean;
  signal ptr_deref_164_store_0_ack_0 : boolean;
  signal ptr_deref_164_store_0_req_1 : boolean;
  signal ptr_deref_164_store_0_ack_1 : boolean;
  signal type_cast_842_inst_ack_1 : boolean;
  signal type_cast_267_inst_ack_1 : boolean;
  signal type_cast_357_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_874_inst_req_1 : boolean;
  signal if_stmt_173_branch_req_0 : boolean;
  signal if_stmt_173_branch_ack_1 : boolean;
  signal if_stmt_173_branch_ack_0 : boolean;
  signal type_cast_198_inst_req_0 : boolean;
  signal type_cast_198_inst_ack_0 : boolean;
  signal type_cast_198_inst_req_1 : boolean;
  signal type_cast_198_inst_ack_1 : boolean;
  signal ptr_deref_467_load_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_856_inst_ack_1 : boolean;
  signal type_cast_185_inst_req_0 : boolean;
  signal array_obj_ref_204_index_offset_req_0 : boolean;
  signal type_cast_947_inst_req_1 : boolean;
  signal array_obj_ref_204_index_offset_ack_0 : boolean;
  signal array_obj_ref_204_index_offset_req_1 : boolean;
  signal array_obj_ref_204_index_offset_ack_1 : boolean;
  signal addr_of_205_final_reg_req_0 : boolean;
  signal addr_of_205_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_874_inst_ack_1 : boolean;
  signal addr_of_205_final_reg_req_1 : boolean;
  signal addr_of_205_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_208_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_208_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_208_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_208_inst_ack_1 : boolean;
  signal type_cast_212_inst_req_0 : boolean;
  signal type_cast_212_inst_ack_0 : boolean;
  signal type_cast_212_inst_req_1 : boolean;
  signal type_cast_212_inst_ack_1 : boolean;
  signal ptr_deref_467_load_0_req_0 : boolean;
  signal type_cast_486_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_856_inst_ack_0 : boolean;
  signal ptr_deref_455_load_0_ack_0 : boolean;
  signal ptr_deref_455_load_0_req_0 : boolean;
  signal type_cast_896_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_856_inst_req_1 : boolean;
  signal ptr_deref_381_load_0_ack_1 : boolean;
  signal ptr_deref_215_store_0_req_0 : boolean;
  signal ptr_deref_215_store_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_910_inst_req_0 : boolean;
  signal ptr_deref_381_load_0_req_1 : boolean;
  signal ptr_deref_215_store_0_req_1 : boolean;
  signal ptr_deref_215_store_0_ack_1 : boolean;
  signal type_cast_486_inst_req_1 : boolean;
  signal type_cast_83_inst_ack_0 : boolean;
  signal ptr_deref_232_load_0_req_0 : boolean;
  signal ptr_deref_232_load_0_ack_0 : boolean;
  signal ptr_deref_232_load_0_req_1 : boolean;
  signal ptr_deref_232_load_0_ack_1 : boolean;
  signal phi_stmt_182_req_0 : boolean;
  signal if_stmt_239_branch_req_0 : boolean;
  signal if_stmt_239_branch_ack_1 : boolean;
  signal if_stmt_239_branch_ack_0 : boolean;
  signal phi_stmt_80_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_249_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_249_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_249_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_249_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_874_inst_req_0 : boolean;
  signal type_cast_253_inst_req_0 : boolean;
  signal type_cast_253_inst_ack_0 : boolean;
  signal type_cast_253_inst_req_1 : boolean;
  signal type_cast_253_inst_ack_1 : boolean;
  signal phi_stmt_150_ack_0 : boolean;
  signal type_cast_896_inst_req_1 : boolean;
  signal ptr_deref_393_load_0_ack_1 : boolean;
  signal ptr_deref_393_load_0_req_1 : boolean;
  signal addr_of_274_final_reg_req_0 : boolean;
  signal addr_of_274_final_reg_ack_0 : boolean;
  signal addr_of_274_final_reg_req_1 : boolean;
  signal addr_of_274_final_reg_ack_1 : boolean;
  signal type_cast_896_inst_ack_1 : boolean;
  signal ptr_deref_277_store_0_ack_0 : boolean;
  signal ptr_deref_381_load_0_req_0 : boolean;
  signal ptr_deref_277_store_0_req_1 : boolean;
  signal ptr_deref_277_store_0_ack_1 : boolean;
  signal ptr_deref_393_load_0_ack_0 : boolean;
  signal ptr_deref_393_load_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_281_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_281_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_281_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_281_inst_ack_1 : boolean;
  signal type_cast_285_inst_req_0 : boolean;
  signal ptr_deref_405_load_0_ack_1 : boolean;
  signal type_cast_285_inst_ack_0 : boolean;
  signal type_cast_285_inst_req_1 : boolean;
  signal type_cast_285_inst_ack_1 : boolean;
  signal type_cast_914_inst_req_1 : boolean;
  signal ptr_deref_368_store_0_ack_1 : boolean;
  signal if_stmt_299_branch_req_0 : boolean;
  signal if_stmt_299_branch_ack_1 : boolean;
  signal if_stmt_299_branch_ack_0 : boolean;
  signal phi_stmt_150_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_910_inst_req_1 : boolean;
  signal type_cast_914_inst_ack_1 : boolean;
  signal STORE_padding_311_store_0_req_0 : boolean;
  signal STORE_padding_311_store_0_ack_0 : boolean;
  signal STORE_padding_311_store_0_req_1 : boolean;
  signal STORE_padding_311_store_0_ack_1 : boolean;
  signal phi_stmt_257_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_315_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_315_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_315_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_315_inst_ack_1 : boolean;
  signal type_cast_319_inst_req_0 : boolean;
  signal type_cast_319_inst_ack_0 : boolean;
  signal type_cast_319_inst_req_1 : boolean;
  signal type_cast_319_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_910_inst_ack_1 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal ptr_deref_330_store_0_req_0 : boolean;
  signal ptr_deref_330_store_0_ack_0 : boolean;
  signal ptr_deref_330_store_0_req_1 : boolean;
  signal ptr_deref_330_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_334_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_334_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_334_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_334_inst_ack_1 : boolean;
  signal type_cast_338_inst_req_0 : boolean;
  signal type_cast_338_inst_ack_0 : boolean;
  signal type_cast_338_inst_req_1 : boolean;
  signal type_cast_338_inst_ack_1 : boolean;
  signal ptr_deref_349_store_0_req_0 : boolean;
  signal ptr_deref_349_store_0_ack_0 : boolean;
  signal ptr_deref_349_store_0_req_1 : boolean;
  signal ptr_deref_349_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_353_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_353_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_353_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_353_inst_ack_1 : boolean;
  signal if_stmt_521_branch_req_0 : boolean;
  signal if_stmt_521_branch_ack_1 : boolean;
  signal if_stmt_521_branch_ack_0 : boolean;
  signal type_cast_540_inst_req_0 : boolean;
  signal type_cast_540_inst_ack_0 : boolean;
  signal type_cast_540_inst_req_1 : boolean;
  signal type_cast_540_inst_ack_1 : boolean;
  signal type_cast_185_inst_ack_1 : boolean;
  signal type_cast_860_inst_ack_1 : boolean;
  signal if_stmt_936_branch_req_0 : boolean;
  signal array_obj_ref_575_index_offset_req_0 : boolean;
  signal array_obj_ref_575_index_offset_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_892_inst_ack_1 : boolean;
  signal array_obj_ref_575_index_offset_req_1 : boolean;
  signal array_obj_ref_575_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_892_inst_req_1 : boolean;
  signal addr_of_576_final_reg_req_0 : boolean;
  signal addr_of_576_final_reg_ack_0 : boolean;
  signal addr_of_576_final_reg_req_1 : boolean;
  signal addr_of_576_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_579_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_579_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_579_inst_req_1 : boolean;
  signal phi_stmt_143_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_579_inst_ack_1 : boolean;
  signal phi_stmt_150_req_1 : boolean;
  signal ptr_deref_922_store_0_ack_1 : boolean;
  signal type_cast_583_inst_req_0 : boolean;
  signal type_cast_583_inst_ack_0 : boolean;
  signal type_cast_583_inst_req_1 : boolean;
  signal type_cast_583_inst_ack_1 : boolean;
  signal type_cast_267_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_892_inst_ack_0 : boolean;
  signal type_cast_263_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_592_inst_req_0 : boolean;
  signal phi_stmt_143_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_592_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_892_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_592_inst_req_1 : boolean;
  signal type_cast_146_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_592_inst_ack_1 : boolean;
  signal ptr_deref_922_store_0_req_1 : boolean;
  signal type_cast_155_inst_ack_1 : boolean;
  signal type_cast_596_inst_req_0 : boolean;
  signal type_cast_146_inst_req_1 : boolean;
  signal type_cast_596_inst_ack_0 : boolean;
  signal type_cast_596_inst_req_1 : boolean;
  signal type_cast_596_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_610_inst_req_0 : boolean;
  signal type_cast_146_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_610_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_610_inst_req_1 : boolean;
  signal type_cast_146_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_610_inst_ack_1 : boolean;
  signal type_cast_263_inst_ack_1 : boolean;
  signal type_cast_155_inst_req_1 : boolean;
  signal type_cast_614_inst_req_0 : boolean;
  signal type_cast_614_inst_ack_0 : boolean;
  signal type_cast_614_inst_req_1 : boolean;
  signal type_cast_614_inst_ack_1 : boolean;
  signal type_cast_267_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_628_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_628_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_628_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_628_inst_ack_1 : boolean;
  signal type_cast_632_inst_req_0 : boolean;
  signal type_cast_632_inst_ack_0 : boolean;
  signal type_cast_632_inst_req_1 : boolean;
  signal type_cast_632_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_646_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_646_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_646_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_646_inst_ack_1 : boolean;
  signal type_cast_263_inst_ack_0 : boolean;
  signal type_cast_155_inst_ack_0 : boolean;
  signal ptr_deref_922_store_0_ack_0 : boolean;
  signal type_cast_650_inst_req_0 : boolean;
  signal type_cast_650_inst_ack_0 : boolean;
  signal type_cast_650_inst_req_1 : boolean;
  signal type_cast_650_inst_ack_1 : boolean;
  signal type_cast_155_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_664_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_664_inst_ack_0 : boolean;
  signal type_cast_878_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_664_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_664_inst_ack_1 : boolean;
  signal type_cast_263_inst_req_0 : boolean;
  signal ptr_deref_922_store_0_req_0 : boolean;
  signal type_cast_668_inst_req_0 : boolean;
  signal type_cast_668_inst_ack_0 : boolean;
  signal type_cast_668_inst_req_1 : boolean;
  signal type_cast_668_inst_ack_1 : boolean;
  signal type_cast_878_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_682_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_682_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_682_inst_req_1 : boolean;
  signal phi_stmt_80_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_682_inst_ack_1 : boolean;
  signal phi_stmt_182_ack_0 : boolean;
  signal type_cast_686_inst_req_0 : boolean;
  signal phi_stmt_73_ack_0 : boolean;
  signal type_cast_686_inst_ack_0 : boolean;
  signal type_cast_686_inst_req_1 : boolean;
  signal type_cast_686_inst_ack_1 : boolean;
  signal phi_stmt_257_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_700_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_700_inst_ack_0 : boolean;
  signal type_cast_878_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_700_inst_req_1 : boolean;
  signal phi_stmt_80_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_700_inst_ack_1 : boolean;
  signal type_cast_185_inst_req_1 : boolean;
  signal type_cast_704_inst_req_0 : boolean;
  signal type_cast_85_inst_ack_1 : boolean;
  signal type_cast_704_inst_ack_0 : boolean;
  signal type_cast_704_inst_req_1 : boolean;
  signal type_cast_85_inst_req_1 : boolean;
  signal type_cast_704_inst_ack_1 : boolean;
  signal type_cast_85_inst_ack_0 : boolean;
  signal type_cast_85_inst_req_0 : boolean;
  signal ptr_deref_712_store_0_req_0 : boolean;
  signal ptr_deref_712_store_0_ack_0 : boolean;
  signal type_cast_860_inst_req_1 : boolean;
  signal ptr_deref_712_store_0_req_1 : boolean;
  signal ptr_deref_712_store_0_ack_1 : boolean;
  signal type_cast_878_inst_req_0 : boolean;
  signal type_cast_185_inst_ack_0 : boolean;
  signal phi_stmt_73_req_0 : boolean;
  signal if_stmt_726_branch_req_0 : boolean;
  signal type_cast_76_inst_ack_1 : boolean;
  signal type_cast_860_inst_ack_0 : boolean;
  signal if_stmt_726_branch_ack_1 : boolean;
  signal type_cast_76_inst_req_1 : boolean;
  signal type_cast_860_inst_req_0 : boolean;
  signal if_stmt_726_branch_ack_0 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal type_cast_750_inst_req_0 : boolean;
  signal type_cast_750_inst_ack_0 : boolean;
  signal type_cast_842_inst_req_1 : boolean;
  signal type_cast_750_inst_req_1 : boolean;
  signal type_cast_750_inst_ack_1 : boolean;
  signal array_obj_ref_785_index_offset_req_0 : boolean;
  signal array_obj_ref_785_index_offset_ack_0 : boolean;
  signal array_obj_ref_785_index_offset_req_1 : boolean;
  signal array_obj_ref_785_index_offset_ack_1 : boolean;
  signal addr_of_786_final_reg_req_0 : boolean;
  signal addr_of_786_final_reg_ack_0 : boolean;
  signal phi_stmt_182_req_1 : boolean;
  signal addr_of_786_final_reg_req_1 : boolean;
  signal addr_of_786_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_789_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_789_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_789_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_789_inst_ack_1 : boolean;
  signal type_cast_793_inst_req_0 : boolean;
  signal type_cast_793_inst_ack_0 : boolean;
  signal type_cast_793_inst_req_1 : boolean;
  signal type_cast_793_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_802_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_802_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_802_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_802_inst_ack_1 : boolean;
  signal type_cast_806_inst_req_0 : boolean;
  signal type_cast_806_inst_ack_0 : boolean;
  signal type_cast_806_inst_req_1 : boolean;
  signal type_cast_806_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_820_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_820_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_820_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_820_inst_ack_1 : boolean;
  signal type_cast_824_inst_req_0 : boolean;
  signal type_cast_824_inst_ack_0 : boolean;
  signal type_cast_824_inst_req_1 : boolean;
  signal type_cast_824_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_838_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_838_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_838_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_838_inst_ack_1 : boolean;
  signal type_cast_842_inst_req_0 : boolean;
  signal type_cast_842_inst_ack_0 : boolean;
  signal type_cast_269_inst_req_0 : boolean;
  signal type_cast_269_inst_ack_0 : boolean;
  signal type_cast_269_inst_req_1 : boolean;
  signal type_cast_269_inst_ack_1 : boolean;
  signal phi_stmt_264_req_1 : boolean;
  signal phi_stmt_257_ack_0 : boolean;
  signal phi_stmt_264_ack_0 : boolean;
  signal type_cast_309_inst_req_0 : boolean;
  signal type_cast_309_inst_ack_0 : boolean;
  signal type_cast_309_inst_req_1 : boolean;
  signal type_cast_309_inst_ack_1 : boolean;
  signal phi_stmt_306_req_0 : boolean;
  signal phi_stmt_306_ack_0 : boolean;
  signal phi_stmt_563_req_0 : boolean;
  signal type_cast_569_inst_req_0 : boolean;
  signal type_cast_569_inst_ack_0 : boolean;
  signal type_cast_569_inst_req_1 : boolean;
  signal type_cast_569_inst_ack_1 : boolean;
  signal phi_stmt_563_req_1 : boolean;
  signal phi_stmt_563_ack_0 : boolean;
  signal phi_stmt_773_req_0 : boolean;
  signal type_cast_779_inst_req_0 : boolean;
  signal type_cast_779_inst_ack_0 : boolean;
  signal type_cast_779_inst_req_1 : boolean;
  signal type_cast_779_inst_ack_1 : boolean;
  signal phi_stmt_773_req_1 : boolean;
  signal phi_stmt_773_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_0: Block -- control-path 
    signal testConfigure_CP_0_elements: BooleanArray(282 downto 0);
    -- 
  begin -- 
    testConfigure_CP_0_elements(0) <= testConfigure_CP_0_start;
    testConfigure_CP_0_symbol <= testConfigure_CP_0_elements(213);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	11 
    -- CP-element group 0:  members (35) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_32/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/branch_block_stmt_32__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/cr
      -- 
    rr_100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_0); -- 
    cr_119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_38_inst_req_1); -- 
    cr_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => ptr_deref_47_store_0_req_1); -- 
    cr_197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_62_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_update_start_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/cr
      -- 
    ra_101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_0, ack => testConfigure_CP_0_elements(1)); -- 
    cr_105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(1), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/rr
      -- 
    ca_106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_1, ack => testConfigure_CP_0_elements(2)); -- 
    rr_114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => type_cast_38_inst_req_0); -- 
    rr_178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => RPIPE_ConvTranspose_input_pipe_58_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/ra
      -- 
    ra_115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_0, ack => testConfigure_CP_0_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/ca
      -- 
    ca_120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_1, ack => testConfigure_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (9) 
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/$exit
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/split_req
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/split_ack
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/rr
      -- 
    rr_158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(5), ack => ptr_deref_47_store_0_req_0); -- 
    testConfigure_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(0) & testConfigure_CP_0_elements(4);
      gj_testConfigure_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/ra
      -- 
    ra_159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_47_store_0_ack_0, ack => testConfigure_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/ca
      -- 
    ca_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_47_store_0_ack_1, ack => testConfigure_CP_0_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_update_start_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/cr
      -- 
    ra_179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_58_inst_ack_0, ack => testConfigure_CP_0_elements(8)); -- 
    cr_183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(8), ack => RPIPE_ConvTranspose_input_pipe_58_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/rr
      -- 
    ca_184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_58_inst_ack_1, ack => testConfigure_CP_0_elements(9)); -- 
    rr_192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(9), ack => type_cast_62_inst_req_0); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/ra
      -- 
    ra_193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_62_inst_ack_0, ack => testConfigure_CP_0_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/ca
      -- 
    ca_198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_62_inst_ack_1, ack => testConfigure_CP_0_elements(11)); -- 
    -- CP-element group 12:  branch  join  transition  place  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	7 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (10) 
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63__exit__
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64__entry__
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_dead_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_eval_test/$entry
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_eval_test/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_eval_test/branch_req
      -- CP-element group 12: 	 branch_block_stmt_32/R_cmp203_65_place
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_if_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_else_link/$entry
      -- 
    branch_req_206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(12), ack => if_stmt_64_branch_req_0); -- 
    testConfigure_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(7) & testConfigure_CP_0_elements(11);
      gj_testConfigure_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  fork  transition  place  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	234 
    -- CP-element group 13: 	235 
    -- CP-element group 13:  members (12) 
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/if_stmt_64_if_link/$exit
      -- CP-element group 13: 	 branch_block_stmt_32/if_stmt_64_if_link/if_choice_transition
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/cr
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/$entry
      -- 
    if_choice_transition_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_64_branch_ack_1, ack => testConfigure_CP_0_elements(13)); -- 
    rr_2462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => type_cast_153_inst_req_0); -- 
    cr_2467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => type_cast_153_inst_req_1); -- 
    -- CP-element group 14:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	221 
    -- CP-element group 14: 	222 
    -- CP-element group 14: 	223 
    -- CP-element group 14:  members (22) 
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70__exit__
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody
      -- CP-element group 14: 	 branch_block_stmt_32/if_stmt_64_else_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/if_stmt_64_else_link/else_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_32/entry_forx_xbodyx_xpreheader
      -- CP-element group 14: 	 branch_block_stmt_32/entry_forx_xbodyx_xpreheader_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/entry_forx_xbodyx_xpreheader_PhiReq/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiAck/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiAck/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiAck/dummy
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiReqMerge
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/cr
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/$entry
      -- 
    else_choice_transition_215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_64_branch_ack_0, ack => testConfigure_CP_0_elements(14)); -- 
    cr_2400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(14), ack => type_cast_85_inst_req_1); -- 
    rr_2395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(14), ack => type_cast_85_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	229 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Sample/ra
      -- 
    ra_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_0, ack => testConfigure_CP_0_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	229 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	31 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Update/ca
      -- 
    ca_234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_1, ack => testConfigure_CP_0_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	229 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	31 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_sample_complete
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Sample/ack
      -- 
    ack_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_101_index_offset_ack_0, ack => testConfigure_CP_0_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	229 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (11) 
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Update/ack
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_request/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_request/req
      -- 
    ack_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_101_index_offset_ack_1, ack => testConfigure_CP_0_elements(18)); -- 
    req_274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(18), ack => addr_of_102_final_reg_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_request/$exit
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_request/ack
      -- 
    ack_275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_102_final_reg_ack_0, ack => testConfigure_CP_0_elements(19)); -- 
    -- CP-element group 20:  join  fork  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	229 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (28) 
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_complete/ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_word_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_root_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_address_resized
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_addr_resize/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_addr_resize/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_addr_resize/base_resize_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_addr_resize/base_resize_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_plus_offset/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_plus_offset/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_plus_offset/sum_rename_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_plus_offset/sum_rename_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_word_addrgen/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_word_addrgen/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_word_addrgen/root_register_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_word_addrgen/root_register_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/ptr_deref_105_Split/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/ptr_deref_105_Split/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/ptr_deref_105_Split/split_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/ptr_deref_105_Split/split_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/word_access_start/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/word_access_start/word_0/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/word_access_start/word_0/rr
      -- 
    ack_280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_102_final_reg_ack_1, ack => testConfigure_CP_0_elements(20)); -- 
    rr_318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(20), ack => ptr_deref_105_store_0_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	30 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/word_access_start/word_0/ra
      -- 
    ra_319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_105_store_0_ack_0, ack => testConfigure_CP_0_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	229 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	31 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/word_access_complete/word_0/ca
      -- 
    ca_330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_105_store_0_ack_1, ack => testConfigure_CP_0_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	229 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/word_access_start/$entry
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/word_access_start/word_0/$entry
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/word_access_start/word_0/rr
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_sample_start_
      -- 
    rr_363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(23), ack => ptr_deref_122_load_0_req_0); -- 
    testConfigure_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(30) & testConfigure_CP_0_elements(229);
      gj_testConfigure_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/word_access_start/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/word_access_start/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/word_access_start/word_0/ra
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_sample_completed_
      -- 
    ra_364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_122_load_0_ack_0, ack => testConfigure_CP_0_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	229 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	31 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/word_access_complete/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/word_access_complete/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/word_access_complete/word_0/ca
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/ptr_deref_122_Merge/$entry
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/ptr_deref_122_Merge/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/ptr_deref_122_Merge/merge_req
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/ptr_deref_122_Merge/merge_ack
      -- 
    ca_375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_122_load_0_ack_1, ack => testConfigure_CP_0_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	229 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_update_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Update/cr
      -- 
    ra_389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_130_inst_ack_0, ack => testConfigure_CP_0_elements(26)); -- 
    cr_393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(26), ack => RPIPE_ConvTranspose_input_pipe_130_inst_req_1); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Sample/rr
      -- 
    ca_394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_130_inst_ack_1, ack => testConfigure_CP_0_elements(27)); -- 
    rr_402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(27), ack => type_cast_134_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Sample/ra
      -- 
    ra_403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_134_inst_ack_0, ack => testConfigure_CP_0_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	229 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Update/ca
      -- 
    ca_408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_134_inst_ack_1, ack => testConfigure_CP_0_elements(29)); -- 
    -- CP-element group 30:  transition  delay-element  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	21 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	23 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_ptr_deref_122_delay
      -- 
    -- Element group testConfigure_CP_0_elements(30) is a control-delay.
    cp_element_30_delay: control_delay_element  generic map(name => " 30_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(21), ack => testConfigure_CP_0_elements(30), clk => clk, reset =>reset);
    -- CP-element group 31:  branch  join  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	16 
    -- CP-element group 31: 	17 
    -- CP-element group 31: 	22 
    -- CP-element group 31: 	25 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (10) 
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135__exit__
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136__entry__
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/$exit
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136_dead_link/$entry
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136_eval_test/$entry
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136_eval_test/$exit
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136_eval_test/branch_req
      -- CP-element group 31: 	 branch_block_stmt_32/R_cmp_137_place
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136_if_link/$entry
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136_else_link/$entry
      -- 
    branch_req_417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(31), ack => if_stmt_136_branch_req_0); -- 
    testConfigure_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(16) & testConfigure_CP_0_elements(17) & testConfigure_CP_0_elements(22) & testConfigure_CP_0_elements(25) & testConfigure_CP_0_elements(29);
      gj_testConfigure_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  place  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	214 
    -- CP-element group 32: 	215 
    -- CP-element group 32: 	217 
    -- CP-element group 32: 	218 
    -- CP-element group 32:  members (20) 
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/cr
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/if_stmt_136_if_link/$exit
      -- CP-element group 32: 	 branch_block_stmt_32/if_stmt_136_if_link/if_choice_transition
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/cr
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/$entry
      -- 
    if_choice_transition_422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_136_branch_ack_1, ack => testConfigure_CP_0_elements(32)); -- 
    rr_2361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_83_inst_req_0); -- 
    cr_2366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_83_inst_req_1); -- 
    rr_2338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_76_inst_req_0); -- 
    cr_2343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_76_inst_req_1); -- 
    -- CP-element group 33:  fork  transition  place  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	230 
    -- CP-element group 33: 	231 
    -- CP-element group 33:  members (12) 
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_136_else_link/$exit
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_136_else_link/else_choice_transition
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Update/cr
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- 
    else_choice_transition_426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_136_branch_ack_0, ack => testConfigure_CP_0_elements(33)); -- 
    cr_2436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(33), ack => type_cast_146_inst_req_1); -- 
    rr_2431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(33), ack => type_cast_146_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	241 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/word_access_start/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/word_access_start/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/word_access_start/word_0/ra
      -- 
    ra_470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_164_store_0_ack_0, ack => testConfigure_CP_0_elements(34)); -- 
    -- CP-element group 35:  branch  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	241 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (15) 
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172__exit__
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173__entry__
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/word_access_complete/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/word_access_complete/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/word_access_complete/word_0/ca
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173_dead_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173_eval_test/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173_eval_test/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173_eval_test/branch_req
      -- CP-element group 35: 	 branch_block_stmt_32/R_cmp12199_174_place
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173_if_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173_else_link/$entry
      -- 
    ca_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_164_store_0_ack_1, ack => testConfigure_CP_0_elements(35)); -- 
    branch_req_489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(35), ack => if_stmt_173_branch_req_0); -- 
    -- CP-element group 36:  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	248 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_32/if_stmt_173_if_link/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/if_stmt_173_if_link/if_choice_transition
      -- CP-element group 36: 	 branch_block_stmt_32/forx_xend_bbx_xnph197
      -- CP-element group 36: 	 branch_block_stmt_32/forx_xend_bbx_xnph197_PhiReq/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/forx_xend_bbx_xnph197_PhiReq/$entry
      -- 
    if_choice_transition_494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_173_branch_ack_1, ack => testConfigure_CP_0_elements(36)); -- 
    -- CP-element group 37:  merge  transition  place  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	245 
    -- CP-element group 37:  members (14) 
      -- CP-element group 37: 	 branch_block_stmt_32/merge_stmt_179__exit__
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_173_else_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_173_else_link/else_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xend_forx_xbody14x_xpreheader
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xend_forx_xbody14x_xpreheader_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xend_forx_xbody14x_xpreheader_PhiReq/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_182/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/merge_stmt_179_PhiAck/dummy
      -- CP-element group 37: 	 branch_block_stmt_32/merge_stmt_179_PhiAck/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/merge_stmt_179_PhiAck/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/merge_stmt_179_PhiReqMerge
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/$entry
      -- 
    else_choice_transition_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_173_branch_ack_0, ack => testConfigure_CP_0_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	247 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Sample/ra
      -- 
    ra_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_198_inst_ack_0, ack => testConfigure_CP_0_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	247 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	55 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Update/ca
      -- 
    ca_517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_198_inst_ack_1, ack => testConfigure_CP_0_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	247 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	55 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_sample_complete
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Sample/ack
      -- 
    ack_543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_204_index_offset_ack_0, ack => testConfigure_CP_0_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	247 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (11) 
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_offset_calculated
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Update/ack
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_request/$entry
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_request/req
      -- 
    ack_548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_204_index_offset_ack_1, ack => testConfigure_CP_0_elements(41)); -- 
    req_557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(41), ack => addr_of_205_final_reg_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_request/$exit
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_request/ack
      -- 
    ack_558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_205_final_reg_ack_0, ack => testConfigure_CP_0_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	247 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	48 
    -- CP-element group 43:  members (19) 
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_complete/ack
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_word_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_root_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_address_resized
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_addr_resize/$entry
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_addr_resize/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_addr_resize/base_resize_req
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_addr_resize/base_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_plus_offset/$entry
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_plus_offset/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_plus_offset/sum_rename_req
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_plus_offset/sum_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_word_addrgen/$entry
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_word_addrgen/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_word_addrgen/root_register_req
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_word_addrgen/root_register_ack
      -- 
    ack_563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_205_final_reg_ack_1, ack => testConfigure_CP_0_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	247 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (6) 
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_update_start_
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Update/cr
      -- 
    ra_572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_208_inst_ack_0, ack => testConfigure_CP_0_elements(44)); -- 
    cr_576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(44), ack => RPIPE_ConvTranspose_input_pipe_208_inst_req_1); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Sample/rr
      -- 
    ca_577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_208_inst_ack_1, ack => testConfigure_CP_0_elements(45)); -- 
    rr_585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(45), ack => type_cast_212_inst_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Sample/ra
      -- 
    ra_586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_212_inst_ack_0, ack => testConfigure_CP_0_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	247 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Update/ca
      -- 
    ca_591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_212_inst_ack_1, ack => testConfigure_CP_0_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	43 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/ptr_deref_215_Split/$entry
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/ptr_deref_215_Split/$exit
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/ptr_deref_215_Split/split_req
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/ptr_deref_215_Split/split_ack
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/word_access_start/$entry
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/word_access_start/word_0/rr
      -- 
    rr_629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(48), ack => ptr_deref_215_store_0_req_0); -- 
    testConfigure_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(43) & testConfigure_CP_0_elements(47);
      gj_testConfigure_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	54 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/word_access_start/word_0/ra
      -- 
    ra_630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_215_store_0_ack_0, ack => testConfigure_CP_0_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	247 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	55 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/word_access_complete/word_0/ca
      -- 
    ca_641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_215_store_0_ack_1, ack => testConfigure_CP_0_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: 	247 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/word_access_start/word_0/rr
      -- 
    rr_674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(51), ack => ptr_deref_232_load_0_req_0); -- 
    testConfigure_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(54) & testConfigure_CP_0_elements(247);
      gj_testConfigure_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/word_access_start/word_0/ra
      -- 
    ra_675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_232_load_0_ack_0, ack => testConfigure_CP_0_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	247 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/word_access_complete/word_0/ca
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/ptr_deref_232_Merge/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/ptr_deref_232_Merge/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/ptr_deref_232_Merge/merge_req
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/ptr_deref_232_Merge/merge_ack
      -- 
    ca_686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_232_load_0_ack_1, ack => testConfigure_CP_0_elements(53)); -- 
    -- CP-element group 54:  transition  delay-element  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	49 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	51 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_ptr_deref_232_delay
      -- 
    -- Element group testConfigure_CP_0_elements(54) is a control-delay.
    cp_element_54_delay: control_delay_element  generic map(name => " 54_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(49), ack => testConfigure_CP_0_elements(54), clk => clk, reset =>reset);
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	50 
    -- CP-element group 55: 	53 
    -- CP-element group 55: 	39 
    -- CP-element group 55: 	40 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238__exit__
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239__entry__
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_32/R_cmp12_240_place
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239_else_link/$entry
      -- 
    branch_req_700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(55), ack => if_stmt_239_branch_req_0); -- 
    testConfigure_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(50) & testConfigure_CP_0_elements(53) & testConfigure_CP_0_elements(39) & testConfigure_CP_0_elements(40);
      gj_testConfigure_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	242 
    -- CP-element group 56: 	243 
    -- CP-element group 56:  members (12) 
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_32/if_stmt_239_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_32/if_stmt_239_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/$entry
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/$entry
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Update/cr
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Update/$entry
      -- 
    if_choice_transition_705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_239_branch_ack_1, ack => testConfigure_CP_0_elements(56)); -- 
    rr_2531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_185_inst_req_0); -- 
    cr_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_185_inst_req_1); -- 
    -- CP-element group 57:  merge  transition  place  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	248 
    -- CP-element group 57:  members (13) 
      -- CP-element group 57: 	 branch_block_stmt_32/merge_stmt_245_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_32/merge_stmt_245_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_32/merge_stmt_245__exit__
      -- CP-element group 57: 	 branch_block_stmt_32/bbx_xnph197x_xloopexit_bbx_xnph197
      -- CP-element group 57: 	 branch_block_stmt_32/merge_stmt_245_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_32/merge_stmt_245_PhiAck/dummy
      -- CP-element group 57: 	 branch_block_stmt_32/if_stmt_239_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_32/if_stmt_239_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_32/forx_xbody14_bbx_xnph197x_xloopexit
      -- CP-element group 57: 	 branch_block_stmt_32/bbx_xnph197x_xloopexit_bbx_xnph197_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_32/bbx_xnph197x_xloopexit_bbx_xnph197_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_32/forx_xbody14_bbx_xnph197x_xloopexit_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_32/forx_xbody14_bbx_xnph197x_xloopexit_PhiReq/$entry
      -- 
    else_choice_transition_709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_239_branch_ack_0, ack => testConfigure_CP_0_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	248 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_update_start_
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Update/cr
      -- 
    ra_723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_249_inst_ack_0, ack => testConfigure_CP_0_elements(58)); -- 
    cr_727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(58), ack => RPIPE_ConvTranspose_input_pipe_249_inst_req_1); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Sample/rr
      -- 
    ca_728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_249_inst_ack_1, ack => testConfigure_CP_0_elements(59)); -- 
    rr_736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(59), ack => type_cast_253_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Sample/ra
      -- 
    ra_737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_253_inst_ack_0, ack => testConfigure_CP_0_elements(60)); -- 
    -- CP-element group 61:  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	248 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	249 
    -- CP-element group 61: 	250 
    -- CP-element group 61: 	251 
    -- CP-element group 61:  members (17) 
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254__exit__
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Update/cr
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_257/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/$entry
      -- 
    ca_742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_253_inst_ack_1, ack => testConfigure_CP_0_elements(61)); -- 
    cr_2609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(61), ack => type_cast_267_inst_req_1); -- 
    rr_2604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(61), ack => type_cast_267_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	264 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_request/$exit
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_request/ack
      -- 
    ack_779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_274_final_reg_ack_0, ack => testConfigure_CP_0_elements(62)); -- 
    -- CP-element group 63:  join  fork  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	264 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (28) 
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_word_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_root_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_address_resized
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_addr_resize/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_addr_resize/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_addr_resize/base_resize_req
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_addr_resize/base_resize_ack
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_plus_offset/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_plus_offset/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_plus_offset/sum_rename_req
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_plus_offset/sum_rename_ack
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_word_addrgen/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_word_addrgen/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_word_addrgen/root_register_req
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_word_addrgen/root_register_ack
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/ptr_deref_277_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/ptr_deref_277_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/ptr_deref_277_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/ptr_deref_277_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/word_access_start/word_0/rr
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_complete/ack
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_sample_start_
      -- 
    ack_784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_274_final_reg_ack_1, ack => testConfigure_CP_0_elements(63)); -- 
    rr_822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(63), ack => ptr_deref_277_store_0_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/word_access_start/word_0/ra
      -- 
    ra_823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_277_store_0_ack_0, ack => testConfigure_CP_0_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	264 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	70 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/word_access_complete/word_0/ca
      -- 
    ca_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_277_store_0_ack_1, ack => testConfigure_CP_0_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	264 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_update_start_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Update/cr
      -- 
    ra_843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_281_inst_ack_0, ack => testConfigure_CP_0_elements(66)); -- 
    cr_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(66), ack => RPIPE_ConvTranspose_input_pipe_281_inst_req_1); -- 
    -- CP-element group 67:  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Sample/rr
      -- 
    ca_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_281_inst_ack_1, ack => testConfigure_CP_0_elements(67)); -- 
    rr_856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(67), ack => type_cast_285_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Sample/ra
      -- 
    ra_857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_285_inst_ack_0, ack => testConfigure_CP_0_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	264 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Update/ca
      -- 
    ca_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_285_inst_ack_1, ack => testConfigure_CP_0_elements(69)); -- 
    -- CP-element group 70:  branch  join  transition  place  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	65 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (10) 
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298__exit__
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299__entry__
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/$exit
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_32/R_exitcond_300_place
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299_else_link/$entry
      -- 
    branch_req_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(70), ack => if_stmt_299_branch_req_0); -- 
    testConfigure_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(65) & testConfigure_CP_0_elements(69);
      gj_testConfigure_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	265 
    -- CP-element group 71: 	266 
    -- CP-element group 71:  members (12) 
      -- CP-element group 71: 	 branch_block_stmt_32/if_stmt_299_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_32/if_stmt_299_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Update/cr
      -- 
    if_choice_transition_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_299_branch_ack_1, ack => testConfigure_CP_0_elements(71)); -- 
    rr_2689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(71), ack => type_cast_309_inst_req_0); -- 
    cr_2694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(71), ack => type_cast_309_inst_req_1); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	254 
    -- CP-element group 72: 	255 
    -- CP-element group 72: 	257 
    -- CP-element group 72: 	258 
    -- CP-element group 72:  members (20) 
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/if_stmt_299_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_32/if_stmt_299_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Update/cr
      -- 
    else_choice_transition_879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_299_branch_ack_0, ack => testConfigure_CP_0_elements(72)); -- 
    cr_2635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_263_inst_req_1); -- 
    rr_2630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_263_inst_req_0); -- 
    rr_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_269_inst_req_0); -- 
    cr_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_269_inst_req_1); -- 
    -- CP-element group 73:  join  fork  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	268 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: 	75 
    -- CP-element group 73: 	76 
    -- CP-element group 73: 	79 
    -- CP-element group 73: 	80 
    -- CP-element group 73: 	82 
    -- CP-element group 73: 	86 
    -- CP-element group 73: 	87 
    -- CP-element group 73: 	89 
    -- CP-element group 73: 	93 
    -- CP-element group 73: 	94 
    -- CP-element group 73: 	96 
    -- CP-element group 73: 	97 
    -- CP-element group 73: 	98 
    -- CP-element group 73: 	99 
    -- CP-element group 73: 	100 
    -- CP-element group 73: 	101 
    -- CP-element group 73: 	102 
    -- CP-element group 73: 	105 
    -- CP-element group 73: 	106 
    -- CP-element group 73: 	107 
    -- CP-element group 73: 	108 
    -- CP-element group 73: 	109 
    -- CP-element group 73: 	110 
    -- CP-element group 73: 	111 
    -- CP-element group 73: 	112 
    -- CP-element group 73: 	113 
    -- CP-element group 73: 	116 
    -- CP-element group 73:  members (280) 
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/STORE_padding_311_Split/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/STORE_padding_311_Split/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/STORE_padding_311_Split/split_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/STORE_padding_311_Split/split_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/word_access_complete/word_0/cr
      -- 
    cr_916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => STORE_padding_311_store_0_req_1); -- 
    rr_905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => STORE_padding_311_store_0_req_0); -- 
    rr_925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => RPIPE_ConvTranspose_input_pipe_315_inst_req_0); -- 
    cr_944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_319_inst_req_1); -- 
    cr_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_330_store_0_req_1); -- 
    cr_1022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_338_inst_req_1); -- 
    cr_1072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_349_store_0_req_1); -- 
    cr_1100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_357_inst_req_1); -- 
    cr_1150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_368_store_0_req_1); -- 
    cr_1195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_381_load_0_req_1); -- 
    rr_1184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_381_load_0_req_0); -- 
    cr_1245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_393_load_0_req_1); -- 
    rr_1234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_393_load_0_req_0); -- 
    cr_1295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_405_load_0_req_1); -- 
    rr_1284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_405_load_0_req_0); -- 
    cr_1314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_419_inst_req_1); -- 
    cr_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_431_load_0_req_1); -- 
    rr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_431_load_0_req_0); -- 
    cr_1409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_443_load_0_req_1); -- 
    rr_1398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_443_load_0_req_0); -- 
    cr_1459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_455_load_0_req_1); -- 
    rr_1448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_455_load_0_req_0); -- 
    cr_1509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_467_load_0_req_1); -- 
    rr_1498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_467_load_0_req_0); -- 
    cr_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_486_inst_req_1); -- 
    testConfigure_CP_0_elements(73) <= testConfigure_CP_0_elements(268);
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/word_access_start/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/word_access_start/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/word_access_start/word_0/ra
      -- 
    ra_906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_311_store_0_ack_0, ack => testConfigure_CP_0_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	119 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/word_access_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/word_access_complete/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/word_access_complete/word_0/ca
      -- 
    ca_917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_311_store_0_ack_1, ack => testConfigure_CP_0_elements(75)); -- 
    -- CP-element group 76:  transition  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	73 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_update_start_
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Update/cr
      -- 
    ra_926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_315_inst_ack_0, ack => testConfigure_CP_0_elements(76)); -- 
    cr_930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(76), ack => RPIPE_ConvTranspose_input_pipe_315_inst_req_1); -- 
    -- CP-element group 77:  fork  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77: 	83 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Update/ca
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Sample/rr
      -- 
    ca_931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_315_inst_ack_1, ack => testConfigure_CP_0_elements(77)); -- 
    rr_939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_319_inst_req_0); -- 
    rr_1003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => RPIPE_ConvTranspose_input_pipe_334_inst_req_0); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Sample/ra
      -- 
    ra_940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_319_inst_ack_0, ack => testConfigure_CP_0_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	73 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Update/ca
      -- 
    ca_945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_319_inst_ack_1, ack => testConfigure_CP_0_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	73 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (9) 
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/ptr_deref_330_Split/$entry
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/ptr_deref_330_Split/$exit
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/ptr_deref_330_Split/split_req
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/ptr_deref_330_Split/split_ack
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/word_access_start/$entry
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/word_access_start/word_0/$entry
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/word_access_start/word_0/rr
      -- 
    rr_983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(80), ack => ptr_deref_330_store_0_req_0); -- 
    testConfigure_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(73) & testConfigure_CP_0_elements(79);
      gj_testConfigure_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	117 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/word_access_start/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/word_access_start/word_0/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/word_access_start/word_0/ra
      -- 
    ra_984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_330_store_0_ack_0, ack => testConfigure_CP_0_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	73 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	119 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/word_access_complete/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/word_access_complete/word_0/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/word_access_complete/word_0/ca
      -- 
    ca_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_330_store_0_ack_1, ack => testConfigure_CP_0_elements(82)); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	77 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_update_start_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Sample/ra
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Update/cr
      -- 
    ra_1004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_334_inst_ack_0, ack => testConfigure_CP_0_elements(83)); -- 
    cr_1008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(83), ack => RPIPE_ConvTranspose_input_pipe_334_inst_req_1); -- 
    -- CP-element group 84:  fork  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	90 
    -- CP-element group 84:  members (9) 
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Sample/rr
      -- 
    ca_1009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_334_inst_ack_1, ack => testConfigure_CP_0_elements(84)); -- 
    rr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(84), ack => type_cast_338_inst_req_0); -- 
    rr_1081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(84), ack => RPIPE_ConvTranspose_input_pipe_353_inst_req_0); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Sample/ra
      -- 
    ra_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_338_inst_ack_0, ack => testConfigure_CP_0_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	73 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Update/ca
      -- 
    ca_1023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_338_inst_ack_1, ack => testConfigure_CP_0_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	73 
    -- CP-element group 87: 	86 
    -- CP-element group 87: 	117 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/ptr_deref_349_Split/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/ptr_deref_349_Split/$exit
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/ptr_deref_349_Split/split_req
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/ptr_deref_349_Split/split_ack
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/word_access_start/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/word_access_start/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/word_access_start/word_0/rr
      -- 
    rr_1061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(87), ack => ptr_deref_349_store_0_req_0); -- 
    testConfigure_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(73) & testConfigure_CP_0_elements(86) & testConfigure_CP_0_elements(117);
      gj_testConfigure_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	118 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/word_access_start/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/word_access_start/word_0/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/word_access_start/word_0/ra
      -- 
    ra_1062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_349_store_0_ack_0, ack => testConfigure_CP_0_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	73 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	119 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/word_access_complete/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/word_access_complete/word_0/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/word_access_complete/word_0/ca
      -- 
    ca_1073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_349_store_0_ack_1, ack => testConfigure_CP_0_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	84 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_update_start_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Update/cr
      -- 
    ra_1082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_353_inst_ack_0, ack => testConfigure_CP_0_elements(90)); -- 
    cr_1086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(90), ack => RPIPE_ConvTranspose_input_pipe_353_inst_req_1); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_sample_start_
      -- 
    ca_1087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_353_inst_ack_1, ack => testConfigure_CP_0_elements(91)); -- 
    rr_1095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(91), ack => type_cast_357_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Sample/ra
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_sample_completed_
      -- 
    ra_1096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_0, ack => testConfigure_CP_0_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	73 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Update/ca
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_update_completed_
      -- 
    ca_1101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_1, ack => testConfigure_CP_0_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	73 
    -- CP-element group 94: 	93 
    -- CP-element group 94: 	118 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/word_access_start/word_0/rr
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/word_access_start/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/word_access_start/$entry
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/ptr_deref_368_Split/split_ack
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/ptr_deref_368_Split/split_req
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/ptr_deref_368_Split/$exit
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/ptr_deref_368_Split/$entry
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/$entry
      -- 
    rr_1139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(94), ack => ptr_deref_368_store_0_req_0); -- 
    testConfigure_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(73) & testConfigure_CP_0_elements(93) & testConfigure_CP_0_elements(118);
      gj_testConfigure_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/word_access_start/word_0/ra
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/word_access_start/word_0/$exit
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/word_access_start/$exit
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/$exit
      -- 
    ra_1140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_368_store_0_ack_0, ack => testConfigure_CP_0_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	73 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	119 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/word_access_complete/word_0/$exit
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/word_access_complete/$exit
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/word_access_complete/word_0/ca
      -- 
    ca_1151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_368_store_0_ack_1, ack => testConfigure_CP_0_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	73 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/word_access_start/word_0/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/word_access_start/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/word_access_start/word_0/ra
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_sample_completed_
      -- 
    ra_1185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_381_load_0_ack_0, ack => testConfigure_CP_0_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	73 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	103 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/ptr_deref_381_Merge/merge_ack
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/ptr_deref_381_Merge/merge_req
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/ptr_deref_381_Merge/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/ptr_deref_381_Merge/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/word_access_complete/word_0/ca
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/word_access_complete/word_0/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/word_access_complete/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/$exit
      -- 
    ca_1196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_381_load_0_ack_1, ack => testConfigure_CP_0_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	73 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/word_access_start/word_0/ra
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/word_access_start/word_0/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/word_access_start/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/$exit
      -- 
    ra_1235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_393_load_0_ack_0, ack => testConfigure_CP_0_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	73 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/word_access_complete/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/ptr_deref_393_Merge/merge_ack
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/ptr_deref_393_Merge/merge_req
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/ptr_deref_393_Merge/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/ptr_deref_393_Merge/$entry
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/word_access_complete/word_0/ca
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/word_access_complete/word_0/$exit
      -- 
    ca_1246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_393_load_0_ack_1, ack => testConfigure_CP_0_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	73 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/word_access_start/word_0/ra
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/word_access_start/word_0/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/word_access_start/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/$exit
      -- 
    ra_1285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_405_load_0_ack_0, ack => testConfigure_CP_0_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	73 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (9) 
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/word_access_complete/word_0/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/word_access_complete/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/ptr_deref_405_Merge/merge_req
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/ptr_deref_405_Merge/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/ptr_deref_405_Merge/merge_ack
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/ptr_deref_405_Merge/$entry
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/word_access_complete/word_0/ca
      -- 
    ca_1296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_405_load_0_ack_1, ack => testConfigure_CP_0_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	98 
    -- CP-element group 103: 	100 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_sample_start_
      -- 
    rr_1309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(103), ack => type_cast_419_inst_req_0); -- 
    testConfigure_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(98) & testConfigure_CP_0_elements(100) & testConfigure_CP_0_elements(102);
      gj_testConfigure_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_sample_completed_
      -- 
    ra_1310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_419_inst_ack_0, ack => testConfigure_CP_0_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	73 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	119 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_update_completed_
      -- 
    ca_1315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_419_inst_ack_1, ack => testConfigure_CP_0_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	73 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (5) 
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/word_access_start/word_0/ra
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/word_access_start/word_0/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/word_access_start/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/$exit
      -- 
    ra_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_431_load_0_ack_0, ack => testConfigure_CP_0_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	73 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	114 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/ptr_deref_431_Merge/merge_ack
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/ptr_deref_431_Merge/merge_req
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/ptr_deref_431_Merge/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/ptr_deref_431_Merge/$entry
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/word_access_complete/word_0/ca
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/word_access_complete/word_0/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/word_access_complete/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/$exit
      -- 
    ca_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_431_load_0_ack_1, ack => testConfigure_CP_0_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	73 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/word_access_start/word_0/ra
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/word_access_start/word_0/$exit
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/word_access_start/$exit
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/$exit
      -- 
    ra_1399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_443_load_0_ack_0, ack => testConfigure_CP_0_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	73 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	114 
    -- CP-element group 109:  members (9) 
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/ptr_deref_443_Merge/merge_ack
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/ptr_deref_443_Merge/merge_req
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/ptr_deref_443_Merge/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/ptr_deref_443_Merge/$entry
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/word_access_complete/word_0/ca
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/word_access_complete/word_0/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/word_access_complete/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/$exit
      -- 
    ca_1410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_443_load_0_ack_1, ack => testConfigure_CP_0_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	73 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/word_access_start/word_0/ra
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/word_access_start/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/word_access_start/$exit
      -- 
    ra_1449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_455_load_0_ack_0, ack => testConfigure_CP_0_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	73 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/word_access_complete/word_0/ca
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/ptr_deref_455_Merge/merge_ack
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/ptr_deref_455_Merge/merge_req
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/ptr_deref_455_Merge/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/ptr_deref_455_Merge/$entry
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/word_access_complete/word_0/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/word_access_complete/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/$exit
      -- 
    ca_1460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_455_load_0_ack_1, ack => testConfigure_CP_0_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	73 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (5) 
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/word_access_start/$exit
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/word_access_start/word_0/ra
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/word_access_start/word_0/$exit
      -- 
    ra_1499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_467_load_0_ack_0, ack => testConfigure_CP_0_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	73 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (9) 
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/word_access_complete/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/ptr_deref_467_Merge/merge_req
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/word_access_complete/word_0/ca
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/ptr_deref_467_Merge/merge_ack
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/ptr_deref_467_Merge/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/word_access_complete/word_0/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/ptr_deref_467_Merge/$entry
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_update_completed_
      -- 
    ca_1510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_467_load_0_ack_1, ack => testConfigure_CP_0_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	107 
    -- CP-element group 114: 	109 
    -- CP-element group 114: 	111 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_sample_start_
      -- 
    rr_1523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(114), ack => type_cast_486_inst_req_0); -- 
    testConfigure_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(107) & testConfigure_CP_0_elements(109) & testConfigure_CP_0_elements(111) & testConfigure_CP_0_elements(113);
      gj_testConfigure_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Sample/ra
      -- 
    ra_1524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_486_inst_ack_0, ack => testConfigure_CP_0_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	73 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	119 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Update/$exit
      -- 
    ca_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_486_inst_ack_1, ack => testConfigure_CP_0_elements(116)); -- 
    -- CP-element group 117:  transition  delay-element  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	81 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	87 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_ptr_deref_349_delay
      -- 
    -- Element group testConfigure_CP_0_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(81), ack => testConfigure_CP_0_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  transition  delay-element  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	88 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	94 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_ptr_deref_368_delay
      -- 
    -- Element group testConfigure_CP_0_elements(118) is a control-delay.
    cp_element_118_delay: control_delay_element  generic map(name => " 118_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(88), ack => testConfigure_CP_0_elements(118), clk => clk, reset =>reset);
    -- CP-element group 119:  branch  join  transition  place  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	75 
    -- CP-element group 119: 	82 
    -- CP-element group 119: 	89 
    -- CP-element group 119: 	96 
    -- CP-element group 119: 	105 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (10) 
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500_eval_test/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500_eval_test/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500_eval_test/branch_req
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500_dead_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/R_cmp65189_501_place
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500_if_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500_else_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499__exit__
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500__entry__
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/$exit
      -- 
    branch_req_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => if_stmt_500_branch_req_0); -- 
    testConfigure_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(75) & testConfigure_CP_0_elements(82) & testConfigure_CP_0_elements(89) & testConfigure_CP_0_elements(96) & testConfigure_CP_0_elements(105) & testConfigure_CP_0_elements(116);
      gj_testConfigure_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	269 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_32/forx_xend37_forx_xcond119x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_32/if_stmt_500_if_link/if_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_32/if_stmt_500_if_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_32/forx_xend37_forx_xcond119x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_32/forx_xend37_forx_xcond119x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_500_branch_ack_1, ack => testConfigure_CP_0_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	124 
    -- CP-element group 121: 	125 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_32/if_stmt_500_else_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/if_stmt_500_else_link/else_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xend37_bbx_xnph191
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_527__exit__
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560__entry__
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_update_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xend37_bbx_xnph191_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xend37_bbx_xnph191_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_527_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_527_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_527_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_527_PhiAck/dummy
      -- 
    else_choice_transition_1548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_500_branch_ack_0, ack => testConfigure_CP_0_elements(121)); -- 
    rr_1583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(121), ack => type_cast_540_inst_req_0); -- 
    cr_1588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(121), ack => type_cast_540_inst_req_1); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	269 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	282 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_32/if_stmt_521_if_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/if_stmt_521_if_link/if_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond119x_xpreheader_forx_xend180
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond119x_xpreheader_forx_xend180_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond119x_xpreheader_forx_xend180_PhiReq/$exit
      -- 
    if_choice_transition_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_521_branch_ack_1, ack => testConfigure_CP_0_elements(122)); -- 
    -- CP-element group 123:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	269 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	168 
    -- CP-element group 123: 	169 
    -- CP-element group 123:  members (18) 
      -- CP-element group 123: 	 branch_block_stmt_32/merge_stmt_732__exit__
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770__entry__
      -- CP-element group 123: 	 branch_block_stmt_32/if_stmt_521_else_link/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/if_stmt_521_else_link/else_choice_transition
      -- CP-element group 123: 	 branch_block_stmt_32/forx_xcond119x_xpreheader_bbx_xnph
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/$entry
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_update_start_
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Sample/rr
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Update/cr
      -- CP-element group 123: 	 branch_block_stmt_32/forx_xcond119x_xpreheader_bbx_xnph_PhiReq/$entry
      -- CP-element group 123: 	 branch_block_stmt_32/forx_xcond119x_xpreheader_bbx_xnph_PhiReq/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/merge_stmt_732_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_32/merge_stmt_732_PhiAck/$entry
      -- CP-element group 123: 	 branch_block_stmt_32/merge_stmt_732_PhiAck/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/merge_stmt_732_PhiAck/dummy
      -- 
    else_choice_transition_1570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_521_branch_ack_0, ack => testConfigure_CP_0_elements(123)); -- 
    rr_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(123), ack => type_cast_750_inst_req_0); -- 
    cr_1947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(123), ack => type_cast_750_inst_req_1); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Sample/ra
      -- 
    ra_1584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_540_inst_ack_0, ack => testConfigure_CP_0_elements(124)); -- 
    -- CP-element group 125:  transition  place  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	121 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	270 
    -- CP-element group 125:  members (9) 
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560__exit__
      -- CP-element group 125: 	 branch_block_stmt_32/bbx_xnph191_forx_xbody67
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_32/bbx_xnph191_forx_xbody67_PhiReq/$entry
      -- CP-element group 125: 	 branch_block_stmt_32/bbx_xnph191_forx_xbody67_PhiReq/phi_stmt_563/$entry
      -- CP-element group 125: 	 branch_block_stmt_32/bbx_xnph191_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/$entry
      -- 
    ca_1589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_540_inst_ack_1, ack => testConfigure_CP_0_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	275 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	165 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_sample_complete
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Sample/ack
      -- 
    ack_1618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_575_index_offset_ack_0, ack => testConfigure_CP_0_elements(126)); -- 
    -- CP-element group 127:  transition  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	275 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (11) 
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_root_address_calculated
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_offset_calculated
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Update/ack
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_base_plus_offset/$entry
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_base_plus_offset/$exit
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_base_plus_offset/sum_rename_req
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_base_plus_offset/sum_rename_ack
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_request/$entry
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_request/req
      -- 
    ack_1623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_575_index_offset_ack_1, ack => testConfigure_CP_0_elements(127)); -- 
    req_1632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(127), ack => addr_of_576_final_reg_req_0); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_request/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_request/ack
      -- 
    ack_1633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_576_final_reg_ack_0, ack => testConfigure_CP_0_elements(128)); -- 
    -- CP-element group 129:  fork  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	275 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	162 
    -- CP-element group 129:  members (19) 
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_complete/$exit
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_complete/ack
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_address_calculated
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_word_address_calculated
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_root_address_calculated
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_address_resized
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_addr_resize/$entry
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_addr_resize/$exit
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_addr_resize/base_resize_req
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_addr_resize/base_resize_ack
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_plus_offset/$entry
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_plus_offset/$exit
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_plus_offset/sum_rename_req
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_plus_offset/sum_rename_ack
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_word_addrgen/$entry
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_word_addrgen/$exit
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_word_addrgen/root_register_req
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_word_addrgen/root_register_ack
      -- 
    ack_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_576_final_reg_ack_1, ack => testConfigure_CP_0_elements(129)); -- 
    -- CP-element group 130:  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	275 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (6) 
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_update_start_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Sample/ra
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Update/cr
      -- 
    ra_1647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_579_inst_ack_0, ack => testConfigure_CP_0_elements(130)); -- 
    cr_1651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(130), ack => RPIPE_ConvTranspose_input_pipe_579_inst_req_1); -- 
    -- CP-element group 131:  fork  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131: 	134 
    -- CP-element group 131:  members (9) 
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Update/ca
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Sample/rr
      -- 
    ca_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_579_inst_ack_1, ack => testConfigure_CP_0_elements(131)); -- 
    rr_1660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(131), ack => type_cast_583_inst_req_0); -- 
    rr_1674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(131), ack => RPIPE_ConvTranspose_input_pipe_592_inst_req_0); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Sample/ra
      -- 
    ra_1661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_583_inst_ack_0, ack => testConfigure_CP_0_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	275 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	162 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Update/ca
      -- 
    ca_1666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_583_inst_ack_1, ack => testConfigure_CP_0_elements(133)); -- 
    -- CP-element group 134:  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	131 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (6) 
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_update_start_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Sample/ra
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Update/cr
      -- 
    ra_1675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_592_inst_ack_0, ack => testConfigure_CP_0_elements(134)); -- 
    cr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(134), ack => RPIPE_ConvTranspose_input_pipe_592_inst_req_1); -- 
    -- CP-element group 135:  fork  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: 	138 
    -- CP-element group 135:  members (9) 
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Update/ca
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Sample/rr
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Sample/rr
      -- 
    ca_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_592_inst_ack_1, ack => testConfigure_CP_0_elements(135)); -- 
    rr_1688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(135), ack => type_cast_596_inst_req_0); -- 
    rr_1702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(135), ack => RPIPE_ConvTranspose_input_pipe_610_inst_req_0); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Sample/ra
      -- 
    ra_1689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_596_inst_ack_0, ack => testConfigure_CP_0_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	275 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	162 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Update/ca
      -- 
    ca_1694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_596_inst_ack_1, ack => testConfigure_CP_0_elements(137)); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	135 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (6) 
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_update_start_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Update/cr
      -- 
    ra_1703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_610_inst_ack_0, ack => testConfigure_CP_0_elements(138)); -- 
    cr_1707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(138), ack => RPIPE_ConvTranspose_input_pipe_610_inst_req_1); -- 
    -- CP-element group 139:  fork  transition  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139: 	142 
    -- CP-element group 139:  members (9) 
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Sample/rr
      -- 
    ca_1708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_610_inst_ack_1, ack => testConfigure_CP_0_elements(139)); -- 
    rr_1716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(139), ack => type_cast_614_inst_req_0); -- 
    rr_1730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(139), ack => RPIPE_ConvTranspose_input_pipe_628_inst_req_0); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Sample/ra
      -- 
    ra_1717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_614_inst_ack_0, ack => testConfigure_CP_0_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	275 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	162 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Update/ca
      -- 
    ca_1722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_614_inst_ack_1, ack => testConfigure_CP_0_elements(141)); -- 
    -- CP-element group 142:  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	139 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (6) 
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_update_start_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Sample/ra
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Update/cr
      -- 
    ra_1731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_628_inst_ack_0, ack => testConfigure_CP_0_elements(142)); -- 
    cr_1735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(142), ack => RPIPE_ConvTranspose_input_pipe_628_inst_req_1); -- 
    -- CP-element group 143:  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143: 	146 
    -- CP-element group 143:  members (9) 
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Update/ca
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Sample/rr
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Sample/rr
      -- 
    ca_1736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_628_inst_ack_1, ack => testConfigure_CP_0_elements(143)); -- 
    rr_1744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(143), ack => type_cast_632_inst_req_0); -- 
    rr_1758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(143), ack => RPIPE_ConvTranspose_input_pipe_646_inst_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Sample/ra
      -- 
    ra_1745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_632_inst_ack_0, ack => testConfigure_CP_0_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	275 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	162 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Update/ca
      -- 
    ca_1750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_632_inst_ack_1, ack => testConfigure_CP_0_elements(145)); -- 
    -- CP-element group 146:  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	143 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (6) 
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_update_start_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Sample/ra
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Update/cr
      -- 
    ra_1759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_646_inst_ack_0, ack => testConfigure_CP_0_elements(146)); -- 
    cr_1763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(146), ack => RPIPE_ConvTranspose_input_pipe_646_inst_req_1); -- 
    -- CP-element group 147:  fork  transition  input  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147: 	150 
    -- CP-element group 147:  members (9) 
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Update/ca
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Sample/rr
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Sample/rr
      -- 
    ca_1764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_646_inst_ack_1, ack => testConfigure_CP_0_elements(147)); -- 
    rr_1772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(147), ack => type_cast_650_inst_req_0); -- 
    rr_1786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(147), ack => RPIPE_ConvTranspose_input_pipe_664_inst_req_0); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Sample/ra
      -- 
    ra_1773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_650_inst_ack_0, ack => testConfigure_CP_0_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	275 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	162 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Update/ca
      -- 
    ca_1778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_650_inst_ack_1, ack => testConfigure_CP_0_elements(149)); -- 
    -- CP-element group 150:  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	147 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (6) 
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_update_start_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Sample/ra
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Update/cr
      -- 
    ra_1787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_664_inst_ack_0, ack => testConfigure_CP_0_elements(150)); -- 
    cr_1791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(150), ack => RPIPE_ConvTranspose_input_pipe_664_inst_req_1); -- 
    -- CP-element group 151:  fork  transition  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151: 	154 
    -- CP-element group 151:  members (9) 
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Update/ca
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Sample/rr
      -- 
    ca_1792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_664_inst_ack_1, ack => testConfigure_CP_0_elements(151)); -- 
    rr_1800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(151), ack => type_cast_668_inst_req_0); -- 
    rr_1814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(151), ack => RPIPE_ConvTranspose_input_pipe_682_inst_req_0); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Sample/ra
      -- 
    ra_1801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_668_inst_ack_0, ack => testConfigure_CP_0_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	275 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	162 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Update/ca
      -- 
    ca_1806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_668_inst_ack_1, ack => testConfigure_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	151 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (6) 
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_update_start_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Update/cr
      -- 
    ra_1815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_682_inst_ack_0, ack => testConfigure_CP_0_elements(154)); -- 
    cr_1819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(154), ack => RPIPE_ConvTranspose_input_pipe_682_inst_req_1); -- 
    -- CP-element group 155:  fork  transition  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	158 
    -- CP-element group 155:  members (9) 
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Sample/rr
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Sample/rr
      -- 
    ca_1820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_682_inst_ack_1, ack => testConfigure_CP_0_elements(155)); -- 
    rr_1828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(155), ack => type_cast_686_inst_req_0); -- 
    rr_1842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(155), ack => RPIPE_ConvTranspose_input_pipe_700_inst_req_0); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Sample/ra
      -- 
    ra_1829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_686_inst_ack_0, ack => testConfigure_CP_0_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	275 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	162 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Update/ca
      -- 
    ca_1834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_686_inst_ack_1, ack => testConfigure_CP_0_elements(157)); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	155 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_update_start_
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Update/cr
      -- 
    ra_1843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_700_inst_ack_0, ack => testConfigure_CP_0_elements(158)); -- 
    cr_1847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(158), ack => RPIPE_ConvTranspose_input_pipe_700_inst_req_1); -- 
    -- CP-element group 159:  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (6) 
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Sample/rr
      -- 
    ca_1848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_700_inst_ack_1, ack => testConfigure_CP_0_elements(159)); -- 
    rr_1856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(159), ack => type_cast_704_inst_req_0); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Sample/ra
      -- 
    ra_1857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_704_inst_ack_0, ack => testConfigure_CP_0_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	275 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Update/ca
      -- 
    ca_1862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_704_inst_ack_1, ack => testConfigure_CP_0_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	129 
    -- CP-element group 162: 	133 
    -- CP-element group 162: 	137 
    -- CP-element group 162: 	141 
    -- CP-element group 162: 	145 
    -- CP-element group 162: 	149 
    -- CP-element group 162: 	153 
    -- CP-element group 162: 	157 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (9) 
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/ptr_deref_712_Split/$entry
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/ptr_deref_712_Split/$exit
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/ptr_deref_712_Split/split_req
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/ptr_deref_712_Split/split_ack
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/word_access_start/$entry
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/word_access_start/word_0/$entry
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/word_access_start/word_0/rr
      -- 
    rr_1900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(162), ack => ptr_deref_712_store_0_req_0); -- 
    testConfigure_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(129) & testConfigure_CP_0_elements(133) & testConfigure_CP_0_elements(137) & testConfigure_CP_0_elements(141) & testConfigure_CP_0_elements(145) & testConfigure_CP_0_elements(149) & testConfigure_CP_0_elements(153) & testConfigure_CP_0_elements(157) & testConfigure_CP_0_elements(161);
      gj_testConfigure_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/word_access_start/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/word_access_start/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/word_access_start/word_0/ra
      -- 
    ra_1901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_712_store_0_ack_0, ack => testConfigure_CP_0_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	275 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/word_access_complete/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/word_access_complete/word_0/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/word_access_complete/word_0/ca
      -- 
    ca_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_712_store_0_ack_1, ack => testConfigure_CP_0_elements(164)); -- 
    -- CP-element group 165:  branch  join  transition  place  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	126 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (10) 
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725__exit__
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726__entry__
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726_dead_link/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726_eval_test/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726_eval_test/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726_eval_test/branch_req
      -- CP-element group 165: 	 branch_block_stmt_32/R_exitcond11_727_place
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726_if_link/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726_else_link/$entry
      -- 
    branch_req_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(165), ack => if_stmt_726_branch_req_0); -- 
    testConfigure_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(126) & testConfigure_CP_0_elements(164);
      gj_testConfigure_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  merge  transition  place  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	269 
    -- CP-element group 166:  members (13) 
      -- CP-element group 166: 	 branch_block_stmt_32/merge_stmt_506__exit__
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader
      -- CP-element group 166: 	 branch_block_stmt_32/if_stmt_726_if_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_32/if_stmt_726_if_link/if_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody67_forx_xcond119x_xpreheaderx_xloopexit
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody67_forx_xcond119x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody67_forx_xcond119x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 166: 	 branch_block_stmt_32/merge_stmt_506_PhiReqMerge
      -- CP-element group 166: 	 branch_block_stmt_32/merge_stmt_506_PhiAck/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/merge_stmt_506_PhiAck/$exit
      -- CP-element group 166: 	 branch_block_stmt_32/merge_stmt_506_PhiAck/dummy
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_726_branch_ack_1, ack => testConfigure_CP_0_elements(166)); -- 
    -- CP-element group 167:  fork  transition  place  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	271 
    -- CP-element group 167: 	272 
    -- CP-element group 167:  members (12) 
      -- CP-element group 167: 	 branch_block_stmt_32/if_stmt_726_else_link/$exit
      -- CP-element group 167: 	 branch_block_stmt_32/if_stmt_726_else_link/else_choice_transition
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_726_branch_ack_0, ack => testConfigure_CP_0_elements(167)); -- 
    rr_2766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(167), ack => type_cast_569_inst_req_0); -- 
    cr_2771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(167), ack => type_cast_569_inst_req_1); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	123 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Sample/ra
      -- 
    ra_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_0, ack => testConfigure_CP_0_elements(168)); -- 
    -- CP-element group 169:  transition  place  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	123 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	276 
    -- CP-element group 169:  members (9) 
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770__exit__
      -- CP-element group 169: 	 branch_block_stmt_32/bbx_xnph_forx_xbody126
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/$exit
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Update/ca
      -- CP-element group 169: 	 branch_block_stmt_32/bbx_xnph_forx_xbody126_PhiReq/$entry
      -- CP-element group 169: 	 branch_block_stmt_32/bbx_xnph_forx_xbody126_PhiReq/phi_stmt_773/$entry
      -- CP-element group 169: 	 branch_block_stmt_32/bbx_xnph_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/$entry
      -- 
    ca_1948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_1, ack => testConfigure_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	281 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	209 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_sample_complete
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Sample/ack
      -- 
    ack_1977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_785_index_offset_ack_0, ack => testConfigure_CP_0_elements(170)); -- 
    -- CP-element group 171:  transition  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	281 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (11) 
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_root_address_calculated
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_offset_calculated
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Update/ack
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_base_plus_offset/$entry
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_base_plus_offset/$exit
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_base_plus_offset/sum_rename_req
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_base_plus_offset/sum_rename_ack
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_request/$entry
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_request/req
      -- 
    ack_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_785_index_offset_ack_1, ack => testConfigure_CP_0_elements(171)); -- 
    req_1991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(171), ack => addr_of_786_final_reg_req_0); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_request/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_request/ack
      -- 
    ack_1992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_786_final_reg_ack_0, ack => testConfigure_CP_0_elements(172)); -- 
    -- CP-element group 173:  fork  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	281 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	206 
    -- CP-element group 173:  members (19) 
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_word_addrgen/root_register_ack
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_word_addrgen/root_register_req
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_word_addrgen/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_word_addrgen/$entry
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_plus_offset/sum_rename_ack
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_plus_offset/sum_rename_req
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_plus_offset/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_plus_offset/$entry
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_addr_resize/base_resize_ack
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_addr_resize/base_resize_req
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_addr_resize/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_addr_resize/$entry
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_address_resized
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_root_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_word_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_complete/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_complete/ack
      -- 
    ack_1997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_786_final_reg_ack_1, ack => testConfigure_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	281 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (6) 
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_update_start_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Sample/ra
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Update/cr
      -- 
    ra_2006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_789_inst_ack_0, ack => testConfigure_CP_0_elements(174)); -- 
    cr_2010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(174), ack => RPIPE_ConvTranspose_input_pipe_789_inst_req_1); -- 
    -- CP-element group 175:  fork  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175: 	178 
    -- CP-element group 175:  members (9) 
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Update/ca
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Sample/rr
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Sample/rr
      -- 
    ca_2011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_789_inst_ack_1, ack => testConfigure_CP_0_elements(175)); -- 
    rr_2019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(175), ack => type_cast_793_inst_req_0); -- 
    rr_2033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(175), ack => RPIPE_ConvTranspose_input_pipe_802_inst_req_0); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Sample/ra
      -- 
    ra_2020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_0, ack => testConfigure_CP_0_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	281 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	206 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Update/ca
      -- 
    ca_2025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_1, ack => testConfigure_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	175 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (6) 
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_update_start_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Sample/ra
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Update/$entry
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Update/cr
      -- 
    ra_2034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_802_inst_ack_0, ack => testConfigure_CP_0_elements(178)); -- 
    cr_2038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(178), ack => RPIPE_ConvTranspose_input_pipe_802_inst_req_1); -- 
    -- CP-element group 179:  fork  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179: 	182 
    -- CP-element group 179:  members (9) 
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Update/ca
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Sample/rr
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Sample/rr
      -- 
    ca_2039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_802_inst_ack_1, ack => testConfigure_CP_0_elements(179)); -- 
    rr_2047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(179), ack => type_cast_806_inst_req_0); -- 
    rr_2061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(179), ack => RPIPE_ConvTranspose_input_pipe_820_inst_req_0); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Sample/ra
      -- 
    ra_2048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_806_inst_ack_0, ack => testConfigure_CP_0_elements(180)); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	281 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	206 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Update/ca
      -- 
    ca_2053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_806_inst_ack_1, ack => testConfigure_CP_0_elements(181)); -- 
    -- CP-element group 182:  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	179 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (6) 
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_update_start_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Sample/ra
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Update/cr
      -- 
    ra_2062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_820_inst_ack_0, ack => testConfigure_CP_0_elements(182)); -- 
    cr_2066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(182), ack => RPIPE_ConvTranspose_input_pipe_820_inst_req_1); -- 
    -- CP-element group 183:  fork  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183: 	186 
    -- CP-element group 183:  members (9) 
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Update/ca
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Sample/rr
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Sample/rr
      -- 
    ca_2067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_820_inst_ack_1, ack => testConfigure_CP_0_elements(183)); -- 
    rr_2075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(183), ack => type_cast_824_inst_req_0); -- 
    rr_2089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(183), ack => RPIPE_ConvTranspose_input_pipe_838_inst_req_0); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Sample/ra
      -- 
    ra_2076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_824_inst_ack_0, ack => testConfigure_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	281 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	206 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Update/ca
      -- 
    ca_2081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_824_inst_ack_1, ack => testConfigure_CP_0_elements(185)); -- 
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	183 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (6) 
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_update_start_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Sample/ra
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Update/cr
      -- 
    ra_2090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_838_inst_ack_0, ack => testConfigure_CP_0_elements(186)); -- 
    cr_2094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(186), ack => RPIPE_ConvTranspose_input_pipe_838_inst_req_1); -- 
    -- CP-element group 187:  fork  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: 	190 
    -- CP-element group 187:  members (9) 
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Sample/rr
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Update/ca
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Sample/rr
      -- 
    ca_2095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_838_inst_ack_1, ack => testConfigure_CP_0_elements(187)); -- 
    rr_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(187), ack => type_cast_842_inst_req_0); -- 
    rr_2117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(187), ack => RPIPE_ConvTranspose_input_pipe_856_inst_req_0); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Sample/ra
      -- 
    ra_2104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_0, ack => testConfigure_CP_0_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	281 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	206 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Update/ca
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_update_completed_
      -- 
    ca_2109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_1, ack => testConfigure_CP_0_elements(189)); -- 
    -- CP-element group 190:  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	187 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (6) 
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_update_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Sample/ra
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Update/cr
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Sample/$exit
      -- 
    ra_2118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_856_inst_ack_0, ack => testConfigure_CP_0_elements(190)); -- 
    cr_2122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(190), ack => RPIPE_ConvTranspose_input_pipe_856_inst_req_1); -- 
    -- CP-element group 191:  fork  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191: 	194 
    -- CP-element group 191:  members (9) 
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Update/ca
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Sample/rr
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Sample/rr
      -- 
    ca_2123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_856_inst_ack_1, ack => testConfigure_CP_0_elements(191)); -- 
    rr_2131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(191), ack => type_cast_860_inst_req_0); -- 
    rr_2145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(191), ack => RPIPE_ConvTranspose_input_pipe_874_inst_req_0); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Sample/ra
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Sample/$exit
      -- 
    ra_2132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_860_inst_ack_0, ack => testConfigure_CP_0_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	281 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	206 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Update/ca
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Update/$exit
      -- 
    ca_2137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_860_inst_ack_1, ack => testConfigure_CP_0_elements(193)); -- 
    -- CP-element group 194:  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	191 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Sample/ra
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Update/cr
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_update_start_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_sample_completed_
      -- 
    ra_2146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_874_inst_ack_0, ack => testConfigure_CP_0_elements(194)); -- 
    cr_2150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(194), ack => RPIPE_ConvTranspose_input_pipe_874_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195: 	198 
    -- CP-element group 195:  members (9) 
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Update/ca
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Sample/rr
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Sample/rr
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Sample/$entry
      -- 
    ca_2151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_874_inst_ack_1, ack => testConfigure_CP_0_elements(195)); -- 
    rr_2159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(195), ack => type_cast_878_inst_req_0); -- 
    rr_2173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(195), ack => RPIPE_ConvTranspose_input_pipe_892_inst_req_0); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Sample/ra
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Sample/$exit
      -- 
    ra_2160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_878_inst_ack_0, ack => testConfigure_CP_0_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	281 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	206 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Update/ca
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_update_completed_
      -- 
    ca_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_878_inst_ack_1, ack => testConfigure_CP_0_elements(197)); -- 
    -- CP-element group 198:  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	195 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (6) 
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Update/cr
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Update/$entry
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Sample/ra
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_update_start_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_sample_completed_
      -- 
    ra_2174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_892_inst_ack_0, ack => testConfigure_CP_0_elements(198)); -- 
    cr_2178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(198), ack => RPIPE_ConvTranspose_input_pipe_892_inst_req_1); -- 
    -- CP-element group 199:  fork  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: 	202 
    -- CP-element group 199:  members (9) 
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Sample/rr
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Sample/rr
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Update/ca
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_update_completed_
      -- 
    ca_2179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_892_inst_ack_1, ack => testConfigure_CP_0_elements(199)); -- 
    rr_2187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(199), ack => type_cast_896_inst_req_0); -- 
    rr_2201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(199), ack => RPIPE_ConvTranspose_input_pipe_910_inst_req_0); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Sample/ra
      -- 
    ra_2188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_896_inst_ack_0, ack => testConfigure_CP_0_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	281 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	206 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Update/ca
      -- 
    ca_2193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_896_inst_ack_1, ack => testConfigure_CP_0_elements(201)); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	199 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Sample/ra
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_sample_completed_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_update_start_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Update/cr
      -- 
    ra_2202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_910_inst_ack_0, ack => testConfigure_CP_0_elements(202)); -- 
    cr_2206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(202), ack => RPIPE_ConvTranspose_input_pipe_910_inst_req_1); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Sample/rr
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_update_completed_
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Update/ca
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_sample_start_
      -- 
    ca_2207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_910_inst_ack_1, ack => testConfigure_CP_0_elements(203)); -- 
    rr_2215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(203), ack => type_cast_914_inst_req_0); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Sample/ra
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_sample_completed_
      -- 
    ra_2216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_914_inst_ack_0, ack => testConfigure_CP_0_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	281 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Update/ca
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_update_completed_
      -- 
    ca_2221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_914_inst_ack_1, ack => testConfigure_CP_0_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	173 
    -- CP-element group 206: 	177 
    -- CP-element group 206: 	181 
    -- CP-element group 206: 	185 
    -- CP-element group 206: 	189 
    -- CP-element group 206: 	193 
    -- CP-element group 206: 	197 
    -- CP-element group 206: 	201 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (9) 
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/word_access_start/word_0/rr
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/word_access_start/word_0/$entry
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/word_access_start/$entry
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/ptr_deref_922_Split/split_ack
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/ptr_deref_922_Split/split_req
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/ptr_deref_922_Split/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/ptr_deref_922_Split/$entry
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/$entry
      -- 
    rr_2259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(206), ack => ptr_deref_922_store_0_req_0); -- 
    testConfigure_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(173) & testConfigure_CP_0_elements(177) & testConfigure_CP_0_elements(181) & testConfigure_CP_0_elements(185) & testConfigure_CP_0_elements(189) & testConfigure_CP_0_elements(193) & testConfigure_CP_0_elements(197) & testConfigure_CP_0_elements(201) & testConfigure_CP_0_elements(205);
      gj_testConfigure_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_sample_completed_
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/word_access_start/word_0/ra
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/word_access_start/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/word_access_start/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/$exit
      -- 
    ra_2260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_922_store_0_ack_0, ack => testConfigure_CP_0_elements(207)); -- 
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	281 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (5) 
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_update_completed_
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/word_access_complete/word_0/ca
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/word_access_complete/word_0/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/word_access_complete/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/$exit
      -- 
    ca_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_922_store_0_ack_1, ack => testConfigure_CP_0_elements(208)); -- 
    -- CP-element group 209:  branch  join  transition  place  output  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	170 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (10) 
      -- CP-element group 209: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935__exit__
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936__entry__
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936_else_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936_if_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936_eval_test/branch_req
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936_eval_test/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936_eval_test/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936_dead_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/R_exitcond19_937_place
      -- CP-element group 209: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/$exit
      -- 
    branch_req_2279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(209), ack => if_stmt_936_branch_req_0); -- 
    testConfigure_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(170) & testConfigure_CP_0_elements(208);
      gj_testConfigure_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  merge  transition  place  input  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	282 
    -- CP-element group 210:  members (13) 
      -- CP-element group 210: 	 branch_block_stmt_32/if_stmt_936_if_link/if_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_32/merge_stmt_942__exit__
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xend180x_xloopexit_forx_xend180
      -- CP-element group 210: 	 branch_block_stmt_32/if_stmt_936_if_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody126_forx_xend180x_xloopexit
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody126_forx_xend180x_xloopexit_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody126_forx_xend180x_xloopexit_PhiReq/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/merge_stmt_942_PhiReqMerge
      -- CP-element group 210: 	 branch_block_stmt_32/merge_stmt_942_PhiAck/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/merge_stmt_942_PhiAck/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/merge_stmt_942_PhiAck/dummy
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xend180x_xloopexit_forx_xend180_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xend180x_xloopexit_forx_xend180_PhiReq/$exit
      -- 
    if_choice_transition_2284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_936_branch_ack_1, ack => testConfigure_CP_0_elements(210)); -- 
    -- CP-element group 211:  fork  transition  place  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	277 
    -- CP-element group 211: 	278 
    -- CP-element group 211:  members (12) 
      -- CP-element group 211: 	 branch_block_stmt_32/if_stmt_936_else_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_32/if_stmt_936_else_link/else_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_936_branch_ack_0, ack => testConfigure_CP_0_elements(211)); -- 
    rr_2820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(211), ack => type_cast_779_inst_req_0); -- 
    cr_2825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(211), ack => type_cast_779_inst_req_1); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	282 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_948/type_cast_947_Sample/ra
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_948/type_cast_947_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_948/type_cast_947_sample_completed_
      -- 
    ra_2302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_947_inst_ack_0, ack => testConfigure_CP_0_elements(212)); -- 
    -- CP-element group 213:  transition  place  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	282 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (16) 
      -- CP-element group 213: 	 $exit
      -- CP-element group 213: 	 branch_block_stmt_32/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/branch_block_stmt_32__exit__
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_948__exit__
      -- CP-element group 213: 	 branch_block_stmt_32/return__
      -- CP-element group 213: 	 branch_block_stmt_32/merge_stmt_950__exit__
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_948/type_cast_947_Update/ca
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_948/type_cast_947_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_948/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_948/type_cast_947_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/return___PhiReq/$entry
      -- CP-element group 213: 	 branch_block_stmt_32/return___PhiReq/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/merge_stmt_950_PhiReqMerge
      -- CP-element group 213: 	 branch_block_stmt_32/merge_stmt_950_PhiAck/$entry
      -- CP-element group 213: 	 branch_block_stmt_32/merge_stmt_950_PhiAck/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/merge_stmt_950_PhiAck/dummy
      -- 
    ca_2307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_947_inst_ack_1, ack => testConfigure_CP_0_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	32 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (2) 
      -- CP-element group 214: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/$exit
      -- CP-element group 214: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/ra
      -- 
    ra_2339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_0, ack => testConfigure_CP_0_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	32 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (2) 
      -- CP-element group 215: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/ca
      -- CP-element group 215: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/$exit
      -- 
    ca_2344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_1, ack => testConfigure_CP_0_elements(215)); -- 
    -- CP-element group 216:  join  transition  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	220 
    -- CP-element group 216:  members (5) 
      -- CP-element group 216: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_req
      -- 
    phi_stmt_73_req_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_73_req_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(216), ack => phi_stmt_73_req_0); -- 
    testConfigure_cp_element_group_216: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_216"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(214) & testConfigure_CP_0_elements(215);
      gj_testConfigure_cp_element_group_216 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	32 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (2) 
      -- CP-element group 217: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/ra
      -- 
    ra_2362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_0, ack => testConfigure_CP_0_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	32 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (2) 
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/ca
      -- 
    ca_2367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_1, ack => testConfigure_CP_0_elements(218)); -- 
    -- CP-element group 219:  join  transition  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_req
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/$exit
      -- 
    phi_stmt_80_req_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_80_req_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(219), ack => phi_stmt_80_req_0); -- 
    testConfigure_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(217) & testConfigure_CP_0_elements(218);
      gj_testConfigure_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  join  transition  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	216 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	226 
    -- CP-element group 220:  members (1) 
      -- CP-element group 220: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_220: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_220"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(216) & testConfigure_CP_0_elements(219);
      gj_testConfigure_cp_element_group_220 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(220), clk => clk, reset => reset); --
    end block;
    -- CP-element group 221:  transition  output  delay-element  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	14 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	225 
    -- CP-element group 221:  members (4) 
      -- CP-element group 221: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_req
      -- CP-element group 221: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_79_konst_delay_trans
      -- 
    phi_stmt_73_req_2379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_73_req_2379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(221), ack => phi_stmt_73_req_1); -- 
    -- Element group testConfigure_CP_0_elements(221) is a control-delay.
    cp_element_221_delay: control_delay_element  generic map(name => " 221_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(14), ack => testConfigure_CP_0_elements(221), clk => clk, reset =>reset);
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	14 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (2) 
      -- CP-element group 222: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/ra
      -- CP-element group 222: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/$exit
      -- 
    ra_2396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_85_inst_ack_0, ack => testConfigure_CP_0_elements(222)); -- 
    -- CP-element group 223:  transition  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	14 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (2) 
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/ca
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/$exit
      -- 
    ca_2401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_85_inst_ack_1, ack => testConfigure_CP_0_elements(223)); -- 
    -- CP-element group 224:  join  transition  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224:  members (5) 
      -- CP-element group 224: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_req
      -- CP-element group 224: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/$exit
      -- 
    phi_stmt_80_req_2402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_80_req_2402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(224), ack => phi_stmt_80_req_1); -- 
    testConfigure_cp_element_group_224: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_224"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(222) & testConfigure_CP_0_elements(223);
      gj_testConfigure_cp_element_group_224 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(224), clk => clk, reset => reset); --
    end block;
    -- CP-element group 225:  join  transition  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	221 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (1) 
      -- CP-element group 225: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(221) & testConfigure_CP_0_elements(224);
      gj_testConfigure_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  merge  fork  transition  place  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	220 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (2) 
      -- CP-element group 226: 	 branch_block_stmt_32/merge_stmt_72_PhiReqMerge
      -- CP-element group 226: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(226) <= OrReduce(testConfigure_CP_0_elements(220) & testConfigure_CP_0_elements(225));
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (1) 
      -- CP-element group 227: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/phi_stmt_73_ack
      -- 
    phi_stmt_73_ack_2407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_73_ack_0, ack => testConfigure_CP_0_elements(227)); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228:  members (1) 
      -- CP-element group 228: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/phi_stmt_80_ack
      -- 
    phi_stmt_80_ack_2408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_80_ack_0, ack => testConfigure_CP_0_elements(228)); -- 
    -- CP-element group 229:  join  fork  transition  place  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	15 
    -- CP-element group 229: 	16 
    -- CP-element group 229: 	17 
    -- CP-element group 229: 	18 
    -- CP-element group 229: 	20 
    -- CP-element group 229: 	22 
    -- CP-element group 229: 	23 
    -- CP-element group 229: 	25 
    -- CP-element group 229: 	26 
    -- CP-element group 229: 	29 
    -- CP-element group 229:  members (61) 
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_72__exit__
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135__entry__
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_word_addrgen/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_word_addrgen/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_word_addrgen/root_register_req
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_word_addrgen/root_register_ack
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_update_start_
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Sample/rr
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Update/cr
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_update_start_
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_resized_1
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_scaled_1
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_computed_1
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_resize_1/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_resize_1/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_resize_1/index_resize_req
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_resize_1/index_resize_ack
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_scale_1/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_scale_1/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_scale_1/scale_rename_req
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_scale_1/scale_rename_ack
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_update_start
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Sample/req
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Update/req
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_complete/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_complete/req
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_update_start_
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/word_access_complete/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/word_access_complete/word_0/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/word_access_complete/word_0/cr
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_update_start_
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_word_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_root_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_address_resized
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_addr_resize/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_addr_resize/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_addr_resize/base_resize_req
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_addr_resize/base_resize_ack
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_plus_offset/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_plus_offset/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_plus_offset/sum_rename_req
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_plus_offset/sum_rename_ack
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/word_access_complete/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/word_access_complete/word_0/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/word_access_complete/word_0/cr
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Sample/rr
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_update_start_
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Update/cr
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/$exit
      -- 
    rr_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(229), ack => type_cast_95_inst_req_0); -- 
    cr_233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(229), ack => type_cast_95_inst_req_1); -- 
    req_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(229), ack => array_obj_ref_101_index_offset_req_0); -- 
    req_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(229), ack => array_obj_ref_101_index_offset_req_1); -- 
    req_279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(229), ack => addr_of_102_final_reg_req_1); -- 
    cr_329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(229), ack => ptr_deref_105_store_0_req_1); -- 
    cr_374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(229), ack => ptr_deref_122_load_0_req_1); -- 
    rr_388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(229), ack => RPIPE_ConvTranspose_input_pipe_130_inst_req_0); -- 
    cr_407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(229), ack => type_cast_134_inst_req_1); -- 
    testConfigure_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(227) & testConfigure_CP_0_elements(228);
      gj_testConfigure_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	33 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230:  members (2) 
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Sample/ra
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Sample/$exit
      -- 
    ra_2432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_146_inst_ack_0, ack => testConfigure_CP_0_elements(230)); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	33 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (2) 
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Update/ca
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Update/$exit
      -- 
    ca_2437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_146_inst_ack_1, ack => testConfigure_CP_0_elements(231)); -- 
    -- CP-element group 232:  join  transition  place  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (8) 
      -- CP-element group 232: 	 branch_block_stmt_32/merge_stmt_142_PhiReqMerge
      -- CP-element group 232: 	 branch_block_stmt_32/merge_stmt_142_PhiAck/$entry
      -- CP-element group 232: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_req
      -- CP-element group 232: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- 
    phi_stmt_143_req_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_143_req_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(232), ack => phi_stmt_143_req_0); -- 
    testConfigure_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(230) & testConfigure_CP_0_elements(231);
      gj_testConfigure_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	237 
    -- CP-element group 233: 	238 
    -- CP-element group 233:  members (13) 
      -- CP-element group 233: 	 branch_block_stmt_32/merge_stmt_142__exit__
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend
      -- CP-element group 233: 	 branch_block_stmt_32/merge_stmt_142_PhiAck/phi_stmt_143_ack
      -- CP-element group 233: 	 branch_block_stmt_32/merge_stmt_142_PhiAck/$exit
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Update/cr
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Sample/rr
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/$entry
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/$entry
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/$entry
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/$entry
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- 
    phi_stmt_143_ack_2443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_143_ack_0, ack => testConfigure_CP_0_elements(233)); -- 
    cr_2493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(233), ack => type_cast_155_inst_req_1); -- 
    rr_2488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(233), ack => type_cast_155_inst_req_0); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	13 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (2) 
      -- CP-element group 234: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/ra
      -- 
    ra_2463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_153_inst_ack_0, ack => testConfigure_CP_0_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	13 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (2) 
      -- CP-element group 235: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/ca
      -- 
    ca_2468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_153_inst_ack_1, ack => testConfigure_CP_0_elements(235)); -- 
    -- CP-element group 236:  join  transition  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	240 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_req
      -- CP-element group 236: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/$exit
      -- 
    phi_stmt_150_req_2469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_150_req_2469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(236), ack => phi_stmt_150_req_0); -- 
    testConfigure_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(234) & testConfigure_CP_0_elements(235);
      gj_testConfigure_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  transition  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	233 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (2) 
      -- CP-element group 237: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Sample/ra
      -- CP-element group 237: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Sample/$exit
      -- 
    ra_2489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_0, ack => testConfigure_CP_0_elements(237)); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	233 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (2) 
      -- CP-element group 238: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Update/ca
      -- CP-element group 238: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Update/$exit
      -- 
    ca_2494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_1, ack => testConfigure_CP_0_elements(238)); -- 
    -- CP-element group 239:  join  transition  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_req
      -- CP-element group 239: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/$exit
      -- CP-element group 239: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/$exit
      -- CP-element group 239: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/$exit
      -- CP-element group 239: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/$exit
      -- CP-element group 239: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    phi_stmt_150_req_2495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_150_req_2495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(239), ack => phi_stmt_150_req_1); -- 
    testConfigure_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(237) & testConfigure_CP_0_elements(238);
      gj_testConfigure_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  merge  transition  place  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	236 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (2) 
      -- CP-element group 240: 	 branch_block_stmt_32/merge_stmt_149_PhiAck/$entry
      -- CP-element group 240: 	 branch_block_stmt_32/merge_stmt_149_PhiReqMerge
      -- 
    testConfigure_CP_0_elements(240) <= OrReduce(testConfigure_CP_0_elements(236) & testConfigure_CP_0_elements(239));
    -- CP-element group 241:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	34 
    -- CP-element group 241: 	35 
    -- CP-element group 241:  members (35) 
      -- CP-element group 241: 	 branch_block_stmt_32/merge_stmt_149__exit__
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172__entry__
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_update_start_
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_address_calculated
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_word_address_calculated
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_root_address_calculated
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_address_resized
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_addr_resize/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_addr_resize/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_addr_resize/base_resize_req
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_addr_resize/base_resize_ack
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_plus_offset/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_plus_offset/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_plus_offset/sum_rename_req
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_plus_offset/sum_rename_ack
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_word_addrgen/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_word_addrgen/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_word_addrgen/root_register_req
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_word_addrgen/root_register_ack
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/ptr_deref_164_Split/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/ptr_deref_164_Split/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/ptr_deref_164_Split/split_req
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/ptr_deref_164_Split/split_ack
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/word_access_start/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/word_access_start/word_0/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/word_access_start/word_0/rr
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/word_access_complete/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/word_access_complete/word_0/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/word_access_complete/word_0/cr
      -- CP-element group 241: 	 branch_block_stmt_32/merge_stmt_149_PhiAck/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/merge_stmt_149_PhiAck/phi_stmt_150_ack
      -- 
    phi_stmt_150_ack_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_150_ack_0, ack => testConfigure_CP_0_elements(241)); -- 
    rr_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => ptr_deref_164_store_0_req_0); -- 
    cr_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => ptr_deref_164_store_0_req_1); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	56 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (2) 
      -- CP-element group 242: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Sample/ra
      -- 
    ra_2532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_185_inst_ack_0, ack => testConfigure_CP_0_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	56 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (2) 
      -- CP-element group 243: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Update/ca
      -- CP-element group 243: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Update/$exit
      -- 
    ca_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_185_inst_ack_1, ack => testConfigure_CP_0_elements(243)); -- 
    -- CP-element group 244:  join  transition  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	246 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_req
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/$exit
      -- 
    phi_stmt_182_req_2538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_182_req_2538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => phi_stmt_182_req_0); -- 
    testConfigure_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(242) & testConfigure_CP_0_elements(243);
      gj_testConfigure_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  transition  output  delay-element  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	37 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (5) 
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/$exit
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_188_konst_delay_trans
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/$exit
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_req
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_182/$exit
      -- 
    phi_stmt_182_req_2549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_182_req_2549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(245), ack => phi_stmt_182_req_1); -- 
    -- Element group testConfigure_CP_0_elements(245) is a control-delay.
    cp_element_245_delay: control_delay_element  generic map(name => " 245_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(37), ack => testConfigure_CP_0_elements(245), clk => clk, reset =>reset);
    -- CP-element group 246:  merge  transition  place  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	244 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (2) 
      -- CP-element group 246: 	 branch_block_stmt_32/merge_stmt_181_PhiAck/$entry
      -- CP-element group 246: 	 branch_block_stmt_32/merge_stmt_181_PhiReqMerge
      -- 
    testConfigure_CP_0_elements(246) <= OrReduce(testConfigure_CP_0_elements(244) & testConfigure_CP_0_elements(245));
    -- CP-element group 247:  fork  transition  place  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	50 
    -- CP-element group 247: 	51 
    -- CP-element group 247: 	53 
    -- CP-element group 247: 	38 
    -- CP-element group 247: 	39 
    -- CP-element group 247: 	40 
    -- CP-element group 247: 	41 
    -- CP-element group 247: 	43 
    -- CP-element group 247: 	44 
    -- CP-element group 247: 	47 
    -- CP-element group 247:  members (62) 
      -- CP-element group 247: 	 branch_block_stmt_32/merge_stmt_181__exit__
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238__entry__
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_update_start_
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Sample/rr
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Update/cr
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_update_start_
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_resized_1
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_scaled_1
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_computed_1
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_resize_1/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_resize_1/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_resize_1/index_resize_req
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_resize_1/index_resize_ack
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_scale_1/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_scale_1/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_scale_1/scale_rename_req
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_scale_1/scale_rename_ack
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_update_start
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Sample/req
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Update/req
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_complete/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_complete/req
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Sample/rr
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_update_start_
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Update/cr
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_update_start_
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/word_access_complete/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/word_access_complete/word_0/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/word_access_complete/word_0/cr
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_update_start_
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_address_calculated
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_word_address_calculated
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_root_address_calculated
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_address_resized
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_addr_resize/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_addr_resize/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_addr_resize/base_resize_req
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_addr_resize/base_resize_ack
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_plus_offset/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_plus_offset/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_plus_offset/sum_rename_req
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_plus_offset/sum_rename_ack
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_word_addrgen/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_word_addrgen/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_word_addrgen/root_register_req
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_word_addrgen/root_register_ack
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/word_access_complete/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/word_access_complete/word_0/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/word_access_complete/word_0/cr
      -- CP-element group 247: 	 branch_block_stmt_32/merge_stmt_181_PhiAck/phi_stmt_182_ack
      -- CP-element group 247: 	 branch_block_stmt_32/merge_stmt_181_PhiAck/$exit
      -- 
    phi_stmt_182_ack_2554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_182_ack_0, ack => testConfigure_CP_0_elements(247)); -- 
    rr_511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(247), ack => type_cast_198_inst_req_0); -- 
    cr_516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(247), ack => type_cast_198_inst_req_1); -- 
    req_542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(247), ack => array_obj_ref_204_index_offset_req_0); -- 
    req_547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(247), ack => array_obj_ref_204_index_offset_req_1); -- 
    req_562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(247), ack => addr_of_205_final_reg_req_1); -- 
    rr_571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(247), ack => RPIPE_ConvTranspose_input_pipe_208_inst_req_0); -- 
    cr_590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(247), ack => type_cast_212_inst_req_1); -- 
    cr_640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(247), ack => ptr_deref_215_store_0_req_1); -- 
    cr_685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(247), ack => ptr_deref_232_load_0_req_1); -- 
    -- CP-element group 248:  merge  fork  transition  place  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	36 
    -- CP-element group 248: 	57 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	58 
    -- CP-element group 248: 	61 
    -- CP-element group 248:  members (13) 
      -- CP-element group 248: 	 branch_block_stmt_32/merge_stmt_247__exit__
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254__entry__
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/$entry
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Sample/rr
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_update_start_
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Update/$entry
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Update/cr
      -- CP-element group 248: 	 branch_block_stmt_32/merge_stmt_247_PhiAck/dummy
      -- CP-element group 248: 	 branch_block_stmt_32/merge_stmt_247_PhiAck/$exit
      -- CP-element group 248: 	 branch_block_stmt_32/merge_stmt_247_PhiAck/$entry
      -- CP-element group 248: 	 branch_block_stmt_32/merge_stmt_247_PhiReqMerge
      -- 
    rr_722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(248), ack => RPIPE_ConvTranspose_input_pipe_249_inst_req_0); -- 
    cr_741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(248), ack => type_cast_253_inst_req_1); -- 
    testConfigure_CP_0_elements(248) <= OrReduce(testConfigure_CP_0_elements(36) & testConfigure_CP_0_elements(57));
    -- CP-element group 249:  transition  output  delay-element  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	61 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	253 
    -- CP-element group 249:  members (4) 
      -- CP-element group 249: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_261_konst_delay_trans
      -- CP-element group 249: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_req
      -- CP-element group 249: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_257/$exit
      -- 
    phi_stmt_257_req_2588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_257_req_2588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => phi_stmt_257_req_0); -- 
    -- Element group testConfigure_CP_0_elements(249) is a control-delay.
    cp_element_249_delay: control_delay_element  generic map(name => " 249_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(61), ack => testConfigure_CP_0_elements(249), clk => clk, reset =>reset);
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	61 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (2) 
      -- CP-element group 250: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Sample/ra
      -- CP-element group 250: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Sample/$exit
      -- 
    ra_2605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_0, ack => testConfigure_CP_0_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	61 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (2) 
      -- CP-element group 251: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Update/ca
      -- 
    ca_2610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_1, ack => testConfigure_CP_0_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (5) 
      -- CP-element group 252: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_req
      -- CP-element group 252: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/$exit
      -- 
    phi_stmt_264_req_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_264_req_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(252), ack => phi_stmt_264_req_0); -- 
    testConfigure_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(250) & testConfigure_CP_0_elements(251);
      gj_testConfigure_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  join  transition  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	249 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	261 
    -- CP-element group 253:  members (1) 
      -- CP-element group 253: 	 branch_block_stmt_32/bbx_xnph197_forx_xbody28_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(249) & testConfigure_CP_0_elements(252);
      gj_testConfigure_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	72 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (2) 
      -- CP-element group 254: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Sample/ra
      -- CP-element group 254: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Sample/$exit
      -- 
    ra_2631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_263_inst_ack_0, ack => testConfigure_CP_0_elements(254)); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	72 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (2) 
      -- CP-element group 255: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Update/$exit
      -- CP-element group 255: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Update/ca
      -- 
    ca_2636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_263_inst_ack_1, ack => testConfigure_CP_0_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	260 
    -- CP-element group 256:  members (5) 
      -- CP-element group 256: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_req
      -- 
    phi_stmt_257_req_2637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_257_req_2637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(256), ack => phi_stmt_257_req_1); -- 
    testConfigure_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(254) & testConfigure_CP_0_elements(255);
      gj_testConfigure_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	72 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (2) 
      -- CP-element group 257: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Sample/ra
      -- 
    ra_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_0, ack => testConfigure_CP_0_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	72 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (2) 
      -- CP-element group 258: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Update/ca
      -- 
    ca_2659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_1, ack => testConfigure_CP_0_elements(258)); -- 
    -- CP-element group 259:  join  transition  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (5) 
      -- CP-element group 259: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_req
      -- 
    phi_stmt_264_req_2660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_264_req_2660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => phi_stmt_264_req_1); -- 
    testConfigure_cp_element_group_259: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_259"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(257) & testConfigure_CP_0_elements(258);
      gj_testConfigure_cp_element_group_259 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 260:  join  transition  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	256 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (1) 
      -- CP-element group 260: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(256) & testConfigure_CP_0_elements(259);
      gj_testConfigure_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  merge  fork  transition  place  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	253 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (2) 
      -- CP-element group 261: 	 branch_block_stmt_32/merge_stmt_256_PhiReqMerge
      -- CP-element group 261: 	 branch_block_stmt_32/merge_stmt_256_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(261) <= OrReduce(testConfigure_CP_0_elements(253) & testConfigure_CP_0_elements(260));
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (1) 
      -- CP-element group 262: 	 branch_block_stmt_32/merge_stmt_256_PhiAck/phi_stmt_257_ack
      -- 
    phi_stmt_257_ack_2665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_257_ack_0, ack => testConfigure_CP_0_elements(262)); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (1) 
      -- CP-element group 263: 	 branch_block_stmt_32/merge_stmt_256_PhiAck/phi_stmt_264_ack
      -- 
    phi_stmt_264_ack_2666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_264_ack_0, ack => testConfigure_CP_0_elements(263)); -- 
    -- CP-element group 264:  join  fork  transition  place  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	62 
    -- CP-element group 264: 	63 
    -- CP-element group 264: 	65 
    -- CP-element group 264: 	66 
    -- CP-element group 264: 	69 
    -- CP-element group 264:  members (42) 
      -- CP-element group 264: 	 branch_block_stmt_32/merge_stmt_256__exit__
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298__entry__
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_update_start_
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_root_address_calculated
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_offset_calculated
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_resized_0
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_scaled_0
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_computed_0
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_resize_0/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_resize_0/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_resize_0/index_resize_req
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_resize_0/index_resize_ack
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_scale_0/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_scale_0/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_scale_0/scale_rename_req
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_scale_0/scale_rename_ack
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_final_index_sum_regn/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_final_index_sum_regn/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_final_index_sum_regn/req
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_final_index_sum_regn/ack
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_base_plus_offset/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_base_plus_offset/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_base_plus_offset/sum_rename_req
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_base_plus_offset/sum_rename_ack
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_request/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_request/req
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_complete/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_complete/req
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_update_start_
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/word_access_complete/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/word_access_complete/word_0/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/word_access_complete/word_0/cr
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Sample/rr
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_update_start_
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_32/merge_stmt_256_PhiAck/$exit
      -- 
    req_778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(264), ack => addr_of_274_final_reg_req_0); -- 
    req_783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(264), ack => addr_of_274_final_reg_req_1); -- 
    cr_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(264), ack => ptr_deref_277_store_0_req_1); -- 
    rr_842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(264), ack => RPIPE_ConvTranspose_input_pipe_281_inst_req_0); -- 
    cr_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(264), ack => type_cast_285_inst_req_1); -- 
    testConfigure_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(262) & testConfigure_CP_0_elements(263);
      gj_testConfigure_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	71 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (2) 
      -- CP-element group 265: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Sample/ra
      -- 
    ra_2690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_309_inst_ack_0, ack => testConfigure_CP_0_elements(265)); -- 
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	71 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (2) 
      -- CP-element group 266: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Update/ca
      -- 
    ca_2695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_309_inst_ack_1, ack => testConfigure_CP_0_elements(266)); -- 
    -- CP-element group 267:  join  transition  place  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (8) 
      -- CP-element group 267: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_req
      -- CP-element group 267: 	 branch_block_stmt_32/merge_stmt_305_PhiReqMerge
      -- CP-element group 267: 	 branch_block_stmt_32/merge_stmt_305_PhiAck/$entry
      -- 
    phi_stmt_306_req_2696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_306_req_2696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => phi_stmt_306_req_0); -- 
    testConfigure_cp_element_group_267: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_267"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(265) & testConfigure_CP_0_elements(266);
      gj_testConfigure_cp_element_group_267 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 268:  merge  transition  place  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	73 
    -- CP-element group 268:  members (4) 
      -- CP-element group 268: 	 branch_block_stmt_32/merge_stmt_305__exit__
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499__entry__
      -- CP-element group 268: 	 branch_block_stmt_32/merge_stmt_305_PhiAck/$exit
      -- CP-element group 268: 	 branch_block_stmt_32/merge_stmt_305_PhiAck/phi_stmt_306_ack
      -- 
    phi_stmt_306_ack_2701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_306_ack_0, ack => testConfigure_CP_0_elements(268)); -- 
    -- CP-element group 269:  merge  branch  transition  place  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	120 
    -- CP-element group 269: 	166 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	122 
    -- CP-element group 269: 	123 
    -- CP-element group 269:  members (17) 
      -- CP-element group 269: 	 branch_block_stmt_32/assign_stmt_514_to_assign_stmt_520/$entry
      -- CP-element group 269: 	 branch_block_stmt_32/assign_stmt_514_to_assign_stmt_520/$exit
      -- CP-element group 269: 	 branch_block_stmt_32/if_stmt_521_dead_link/$entry
      -- CP-element group 269: 	 branch_block_stmt_32/if_stmt_521_eval_test/$entry
      -- CP-element group 269: 	 branch_block_stmt_32/merge_stmt_508__exit__
      -- CP-element group 269: 	 branch_block_stmt_32/assign_stmt_514_to_assign_stmt_520__entry__
      -- CP-element group 269: 	 branch_block_stmt_32/assign_stmt_514_to_assign_stmt_520__exit__
      -- CP-element group 269: 	 branch_block_stmt_32/if_stmt_521__entry__
      -- CP-element group 269: 	 branch_block_stmt_32/if_stmt_521_eval_test/$exit
      -- CP-element group 269: 	 branch_block_stmt_32/if_stmt_521_eval_test/branch_req
      -- CP-element group 269: 	 branch_block_stmt_32/R_cmp124185_522_place
      -- CP-element group 269: 	 branch_block_stmt_32/if_stmt_521_if_link/$entry
      -- CP-element group 269: 	 branch_block_stmt_32/if_stmt_521_else_link/$entry
      -- CP-element group 269: 	 branch_block_stmt_32/merge_stmt_508_PhiReqMerge
      -- CP-element group 269: 	 branch_block_stmt_32/merge_stmt_508_PhiAck/$entry
      -- CP-element group 269: 	 branch_block_stmt_32/merge_stmt_508_PhiAck/$exit
      -- CP-element group 269: 	 branch_block_stmt_32/merge_stmt_508_PhiAck/dummy
      -- 
    branch_req_1561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(269), ack => if_stmt_521_branch_req_0); -- 
    testConfigure_CP_0_elements(269) <= OrReduce(testConfigure_CP_0_elements(120) & testConfigure_CP_0_elements(166));
    -- CP-element group 270:  transition  output  delay-element  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	125 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	274 
    -- CP-element group 270:  members (5) 
      -- CP-element group 270: 	 branch_block_stmt_32/bbx_xnph191_forx_xbody67_PhiReq/$exit
      -- CP-element group 270: 	 branch_block_stmt_32/bbx_xnph191_forx_xbody67_PhiReq/phi_stmt_563/$exit
      -- CP-element group 270: 	 branch_block_stmt_32/bbx_xnph191_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/$exit
      -- CP-element group 270: 	 branch_block_stmt_32/bbx_xnph191_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_567_konst_delay_trans
      -- CP-element group 270: 	 branch_block_stmt_32/bbx_xnph191_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_req
      -- 
    phi_stmt_563_req_2747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_563_req_2747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(270), ack => phi_stmt_563_req_0); -- 
    -- Element group testConfigure_CP_0_elements(270) is a control-delay.
    cp_element_270_delay: control_delay_element  generic map(name => " 270_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(125), ack => testConfigure_CP_0_elements(270), clk => clk, reset =>reset);
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	167 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	273 
    -- CP-element group 271:  members (2) 
      -- CP-element group 271: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Sample/ra
      -- 
    ra_2767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_569_inst_ack_0, ack => testConfigure_CP_0_elements(271)); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	167 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (2) 
      -- CP-element group 272: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Update/ca
      -- 
    ca_2772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_569_inst_ack_1, ack => testConfigure_CP_0_elements(272)); -- 
    -- CP-element group 273:  join  transition  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	271 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/$exit
      -- CP-element group 273: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/$exit
      -- CP-element group 273: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/$exit
      -- CP-element group 273: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/$exit
      -- CP-element group 273: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/$exit
      -- CP-element group 273: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_req
      -- 
    phi_stmt_563_req_2773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_563_req_2773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(273), ack => phi_stmt_563_req_1); -- 
    testConfigure_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(271) & testConfigure_CP_0_elements(272);
      gj_testConfigure_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  merge  transition  place  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	270 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (2) 
      -- CP-element group 274: 	 branch_block_stmt_32/merge_stmt_562_PhiReqMerge
      -- CP-element group 274: 	 branch_block_stmt_32/merge_stmt_562_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(274) <= OrReduce(testConfigure_CP_0_elements(270) & testConfigure_CP_0_elements(273));
    -- CP-element group 275:  fork  transition  place  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	126 
    -- CP-element group 275: 	127 
    -- CP-element group 275: 	129 
    -- CP-element group 275: 	130 
    -- CP-element group 275: 	133 
    -- CP-element group 275: 	137 
    -- CP-element group 275: 	141 
    -- CP-element group 275: 	145 
    -- CP-element group 275: 	149 
    -- CP-element group 275: 	153 
    -- CP-element group 275: 	157 
    -- CP-element group 275: 	161 
    -- CP-element group 275: 	164 
    -- CP-element group 275:  members (56) 
      -- CP-element group 275: 	 branch_block_stmt_32/merge_stmt_562__exit__
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725__entry__
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_resized_1
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_scaled_1
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_computed_1
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_resize_1/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_resize_1/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_resize_1/index_resize_req
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_resize_1/index_resize_ack
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_scale_1/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_scale_1/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_scale_1/scale_rename_req
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_scale_1/scale_rename_ack
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_update_start
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Sample/req
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Update/req
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_complete/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_complete/req
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Sample/rr
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/word_access_complete/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/word_access_complete/word_0/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/word_access_complete/word_0/cr
      -- CP-element group 275: 	 branch_block_stmt_32/merge_stmt_562_PhiAck/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/merge_stmt_562_PhiAck/phi_stmt_563_ack
      -- 
    phi_stmt_563_ack_2778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_563_ack_0, ack => testConfigure_CP_0_elements(275)); -- 
    req_1617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => array_obj_ref_575_index_offset_req_0); -- 
    req_1622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => array_obj_ref_575_index_offset_req_1); -- 
    req_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => addr_of_576_final_reg_req_1); -- 
    rr_1646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => RPIPE_ConvTranspose_input_pipe_579_inst_req_0); -- 
    cr_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => type_cast_583_inst_req_1); -- 
    cr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => type_cast_596_inst_req_1); -- 
    cr_1721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => type_cast_614_inst_req_1); -- 
    cr_1749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => type_cast_632_inst_req_1); -- 
    cr_1777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => type_cast_650_inst_req_1); -- 
    cr_1805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => type_cast_668_inst_req_1); -- 
    cr_1833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => type_cast_686_inst_req_1); -- 
    cr_1861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => type_cast_704_inst_req_1); -- 
    cr_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => ptr_deref_712_store_0_req_1); -- 
    -- CP-element group 276:  transition  output  delay-element  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	169 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	280 
    -- CP-element group 276:  members (5) 
      -- CP-element group 276: 	 branch_block_stmt_32/bbx_xnph_forx_xbody126_PhiReq/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/bbx_xnph_forx_xbody126_PhiReq/phi_stmt_773/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/bbx_xnph_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/bbx_xnph_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_777_konst_delay_trans
      -- CP-element group 276: 	 branch_block_stmt_32/bbx_xnph_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_req
      -- 
    phi_stmt_773_req_2801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_773_req_2801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(276), ack => phi_stmt_773_req_0); -- 
    -- Element group testConfigure_CP_0_elements(276) is a control-delay.
    cp_element_276_delay: control_delay_element  generic map(name => " 276_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(169), ack => testConfigure_CP_0_elements(276), clk => clk, reset =>reset);
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	211 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (2) 
      -- CP-element group 277: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Sample/ra
      -- 
    ra_2821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_779_inst_ack_0, ack => testConfigure_CP_0_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	211 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (2) 
      -- CP-element group 278: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Update/ca
      -- 
    ca_2826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_779_inst_ack_1, ack => testConfigure_CP_0_elements(278)); -- 
    -- CP-element group 279:  join  transition  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_req
      -- 
    phi_stmt_773_req_2827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_773_req_2827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(279), ack => phi_stmt_773_req_1); -- 
    testConfigure_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(277) & testConfigure_CP_0_elements(278);
      gj_testConfigure_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  merge  transition  place  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	276 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (2) 
      -- CP-element group 280: 	 branch_block_stmt_32/merge_stmt_772_PhiReqMerge
      -- CP-element group 280: 	 branch_block_stmt_32/merge_stmt_772_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(280) <= OrReduce(testConfigure_CP_0_elements(276) & testConfigure_CP_0_elements(279));
    -- CP-element group 281:  fork  transition  place  input  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	170 
    -- CP-element group 281: 	171 
    -- CP-element group 281: 	173 
    -- CP-element group 281: 	174 
    -- CP-element group 281: 	177 
    -- CP-element group 281: 	181 
    -- CP-element group 281: 	185 
    -- CP-element group 281: 	189 
    -- CP-element group 281: 	193 
    -- CP-element group 281: 	197 
    -- CP-element group 281: 	201 
    -- CP-element group 281: 	205 
    -- CP-element group 281: 	208 
    -- CP-element group 281:  members (56) 
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_update_start_
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/merge_stmt_772__exit__
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935__entry__
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Update/cr
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Update/cr
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_update_start_
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_update_start_
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/word_access_complete/word_0/cr
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/word_access_complete/word_0/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/word_access_complete/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Update/cr
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_update_start_
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Update/cr
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Update/cr
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_update_start_
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_resized_1
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_scaled_1
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_computed_1
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_resize_1/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_resize_1/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_resize_1/index_resize_req
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_resize_1/index_resize_ack
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_scale_1/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_scale_1/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_scale_1/scale_rename_req
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_scale_1/scale_rename_ack
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_update_start
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Sample/req
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Update/req
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_update_start_
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_complete/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_complete/req
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_sample_start_
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Sample/rr
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_update_start_
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Update/cr
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_update_start_
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Update/cr
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_update_start_
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Update/cr
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_update_start_
      -- CP-element group 281: 	 branch_block_stmt_32/merge_stmt_772_PhiAck/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/merge_stmt_772_PhiAck/phi_stmt_773_ack
      -- 
    phi_stmt_773_ack_2832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_773_ack_0, ack => testConfigure_CP_0_elements(281)); -- 
    cr_2192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => type_cast_896_inst_req_1); -- 
    cr_2220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => type_cast_914_inst_req_1); -- 
    cr_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => ptr_deref_922_store_0_req_1); -- 
    cr_2164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => type_cast_878_inst_req_1); -- 
    cr_2136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => type_cast_860_inst_req_1); -- 
    cr_2108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => type_cast_842_inst_req_1); -- 
    req_1976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => array_obj_ref_785_index_offset_req_0); -- 
    req_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => array_obj_ref_785_index_offset_req_1); -- 
    req_1996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => addr_of_786_final_reg_req_1); -- 
    rr_2005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => RPIPE_ConvTranspose_input_pipe_789_inst_req_0); -- 
    cr_2024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => type_cast_793_inst_req_1); -- 
    cr_2052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => type_cast_806_inst_req_1); -- 
    cr_2080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => type_cast_824_inst_req_1); -- 
    -- CP-element group 282:  merge  fork  transition  place  output  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	122 
    -- CP-element group 282: 	210 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	212 
    -- CP-element group 282: 	213 
    -- CP-element group 282:  members (13) 
      -- CP-element group 282: 	 branch_block_stmt_32/assign_stmt_948/$entry
      -- CP-element group 282: 	 branch_block_stmt_32/merge_stmt_944__exit__
      -- CP-element group 282: 	 branch_block_stmt_32/assign_stmt_948__entry__
      -- CP-element group 282: 	 branch_block_stmt_32/assign_stmt_948/type_cast_947_Sample/rr
      -- CP-element group 282: 	 branch_block_stmt_32/assign_stmt_948/type_cast_947_sample_start_
      -- CP-element group 282: 	 branch_block_stmt_32/assign_stmt_948/type_cast_947_Sample/$entry
      -- CP-element group 282: 	 branch_block_stmt_32/assign_stmt_948/type_cast_947_Update/$entry
      -- CP-element group 282: 	 branch_block_stmt_32/assign_stmt_948/type_cast_947_Update/cr
      -- CP-element group 282: 	 branch_block_stmt_32/assign_stmt_948/type_cast_947_update_start_
      -- CP-element group 282: 	 branch_block_stmt_32/merge_stmt_944_PhiReqMerge
      -- CP-element group 282: 	 branch_block_stmt_32/merge_stmt_944_PhiAck/$entry
      -- CP-element group 282: 	 branch_block_stmt_32/merge_stmt_944_PhiAck/$exit
      -- CP-element group 282: 	 branch_block_stmt_32/merge_stmt_944_PhiAck/dummy
      -- 
    rr_2301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(282), ack => type_cast_947_inst_req_0); -- 
    cr_2306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(282), ack => type_cast_947_inst_req_1); -- 
    testConfigure_CP_0_elements(282) <= OrReduce(testConfigure_CP_0_elements(122) & testConfigure_CP_0_elements(210));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar215_574_resized : std_logic_vector(13 downto 0);
    signal R_indvar215_574_scaled : std_logic_vector(13 downto 0);
    signal R_indvar225_272_resized : std_logic_vector(0 downto 0);
    signal R_indvar225_272_scaled : std_logic_vector(0 downto 0);
    signal R_indvar228_203_resized : std_logic_vector(6 downto 0);
    signal R_indvar228_203_scaled : std_logic_vector(6 downto 0);
    signal R_indvar233_100_resized : std_logic_vector(6 downto 0);
    signal R_indvar233_100_scaled : std_logic_vector(6 downto 0);
    signal R_indvar_784_resized : std_logic_vector(10 downto 0);
    signal R_indvar_784_scaled : std_logic_vector(10 downto 0);
    signal STORE_padding_311_data_0 : std_logic_vector(15 downto 0);
    signal STORE_padding_311_word_address_0 : std_logic_vector(0 downto 0);
    signal add104_692 : std_logic_vector(63 downto 0);
    signal add110_710 : std_logic_vector(63 downto 0);
    signal add136_812 : std_logic_vector(63 downto 0);
    signal add142_830 : std_logic_vector(63 downto 0);
    signal add148_848 : std_logic_vector(63 downto 0);
    signal add154_866 : std_logic_vector(63 downto 0);
    signal add160_884 : std_logic_vector(63 downto 0);
    signal add166_902 : std_logic_vector(63 downto 0);
    signal add172_920 : std_logic_vector(63 downto 0);
    signal add80_620 : std_logic_vector(63 downto 0);
    signal add86_638 : std_logic_vector(63 downto 0);
    signal add92_656 : std_logic_vector(63 downto 0);
    signal add98_674 : std_logic_vector(63 downto 0);
    signal add_602 : std_logic_vector(63 downto 0);
    signal array_obj_ref_101_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_204_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_204_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_204_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_204_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_204_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_204_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_273_final_offset : std_logic_vector(0 downto 0);
    signal array_obj_ref_273_offset_scale_factor_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_273_resized_base_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_273_root_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_575_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_575_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_575_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_575_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_575_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_575_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_785_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_785_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_785_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_785_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_785_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_785_root_address : std_logic_vector(10 downto 0);
    signal arrayidx114_577 : std_logic_vector(31 downto 0);
    signal arrayidx176_787 : std_logic_vector(31 downto 0);
    signal arrayidx19_206 : std_logic_vector(31 downto 0);
    signal arrayidx33_275 : std_logic_vector(31 downto 0);
    signal arrayidx_103 : std_logic_vector(31 downto 0);
    signal call101_683 : std_logic_vector(7 downto 0);
    signal call107_701 : std_logic_vector(7 downto 0);
    signal call129_790 : std_logic_vector(7 downto 0);
    signal call133_803 : std_logic_vector(7 downto 0);
    signal call139_821 : std_logic_vector(7 downto 0);
    signal call145_839 : std_logic_vector(7 downto 0);
    signal call151_857 : std_logic_vector(7 downto 0);
    signal call157_875 : std_logic_vector(7 downto 0);
    signal call15_209 : std_logic_vector(7 downto 0);
    signal call163_893 : std_logic_vector(7 downto 0);
    signal call169_911 : std_logic_vector(7 downto 0);
    signal call29193_250 : std_logic_vector(7 downto 0);
    signal call29_282 : std_logic_vector(7 downto 0);
    signal call3204_59 : std_logic_vector(7 downto 0);
    signal call3_131 : std_logic_vector(7 downto 0);
    signal call40_316 : std_logic_vector(7 downto 0);
    signal call42_335 : std_logic_vector(7 downto 0);
    signal call44_354 : std_logic_vector(7 downto 0);
    signal call69_580 : std_logic_vector(7 downto 0);
    signal call72_593 : std_logic_vector(7 downto 0);
    signal call77_611 : std_logic_vector(7 downto 0);
    signal call83_629 : std_logic_vector(7 downto 0);
    signal call89_647 : std_logic_vector(7 downto 0);
    signal call95_665 : std_logic_vector(7 downto 0);
    signal call_35 : std_logic_vector(7 downto 0);
    signal cmp12199_172 : std_logic_vector(0 downto 0);
    signal cmp124185_520 : std_logic_vector(0 downto 0);
    signal cmp12_238 : std_logic_vector(0 downto 0);
    signal cmp203_56 : std_logic_vector(0 downto 0);
    signal cmp65189_499 : std_logic_vector(0 downto 0);
    signal cmp_128 : std_logic_vector(0 downto 0);
    signal conv103_687 : std_logic_vector(63 downto 0);
    signal conv109_705 : std_logic_vector(63 downto 0);
    signal conv130_794 : std_logic_vector(63 downto 0);
    signal conv135_807 : std_logic_vector(63 downto 0);
    signal conv141_825 : std_logic_vector(63 downto 0);
    signal conv147_843 : std_logic_vector(63 downto 0);
    signal conv153_861 : std_logic_vector(63 downto 0);
    signal conv159_879 : std_logic_vector(63 downto 0);
    signal conv165_897 : std_logic_vector(63 downto 0);
    signal conv16_213 : std_logic_vector(31 downto 0);
    signal conv171_915 : std_logic_vector(63 downto 0);
    signal conv30194_254 : std_logic_vector(15 downto 0);
    signal conv30196_264 : std_logic_vector(15 downto 0);
    signal conv30_286 : std_logic_vector(15 downto 0);
    signal conv30x_xlcssa_306 : std_logic_vector(15 downto 0);
    signal conv41_320 : std_logic_vector(31 downto 0);
    signal conv4205_63 : std_logic_vector(31 downto 0);
    signal conv4207_80 : std_logic_vector(31 downto 0);
    signal conv43_339 : std_logic_vector(31 downto 0);
    signal conv45_358 : std_logic_vector(31 downto 0);
    signal conv4_135 : std_logic_vector(31 downto 0);
    signal conv4x_xlcssa1_143 : std_logic_vector(31 downto 0);
    signal conv4x_xlcssa_150 : std_logic_vector(31 downto 0);
    signal conv51_420 : std_logic_vector(63 downto 0);
    signal conv60_487 : std_logic_vector(63 downto 0);
    signal conv70_584 : std_logic_vector(63 downto 0);
    signal conv74_597 : std_logic_vector(63 downto 0);
    signal conv79_615 : std_logic_vector(63 downto 0);
    signal conv85_633 : std_logic_vector(63 downto 0);
    signal conv91_651 : std_logic_vector(63 downto 0);
    signal conv97_669 : std_logic_vector(63 downto 0);
    signal conv_39 : std_logic_vector(31 downto 0);
    signal exitcond11_725 : std_logic_vector(0 downto 0);
    signal exitcond19_935 : std_logic_vector(0 downto 0);
    signal exitcond_298 : std_logic_vector(0 downto 0);
    signal iNsTr_13_119 : std_logic_vector(31 downto 0);
    signal iNsTr_1_45 : std_logic_vector(31 downto 0);
    signal iNsTr_21_229 : std_logic_vector(31 downto 0);
    signal iNsTr_26_328 : std_logic_vector(31 downto 0);
    signal iNsTr_29_347 : std_logic_vector(31 downto 0);
    signal iNsTr_32_366 : std_logic_vector(31 downto 0);
    signal iNsTr_34_378 : std_logic_vector(31 downto 0);
    signal iNsTr_35_390 : std_logic_vector(31 downto 0);
    signal iNsTr_36_402 : std_logic_vector(31 downto 0);
    signal iNsTr_37_428 : std_logic_vector(31 downto 0);
    signal iNsTr_38_440 : std_logic_vector(31 downto 0);
    signal iNsTr_39_452 : std_logic_vector(31 downto 0);
    signal iNsTr_40_464 : std_logic_vector(31 downto 0);
    signal iNsTr_5_162 : std_logic_vector(31 downto 0);
    signal inc22_199 : std_logic_vector(31 downto 0);
    signal inc_96 : std_logic_vector(31 downto 0);
    signal indvar215_563 : std_logic_vector(63 downto 0);
    signal indvar225_257 : std_logic_vector(63 downto 0);
    signal indvar228_182 : std_logic_vector(63 downto 0);
    signal indvar233_73 : std_logic_vector(63 downto 0);
    signal indvar_773 : std_logic_vector(63 downto 0);
    signal indvarx_xnext216_720 : std_logic_vector(63 downto 0);
    signal indvarx_xnext226_292 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_930 : std_logic_vector(63 downto 0);
    signal mul50_416 : std_logic_vector(31 downto 0);
    signal mul55_473 : std_logic_vector(31 downto 0);
    signal mul57_478 : std_logic_vector(31 downto 0);
    signal mul59_483 : std_logic_vector(31 downto 0);
    signal mul_411 : std_logic_vector(31 downto 0);
    signal ptr_deref_105_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_105_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_105_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_105_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_105_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_105_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_122_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_122_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_122_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_122_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_122_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_164_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_164_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_164_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_164_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_164_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_164_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_215_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_215_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_215_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_215_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_215_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_215_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_232_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_232_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_232_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_232_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_232_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_277_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_277_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_277_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_277_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_277_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_277_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_330_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_330_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_330_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_330_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_330_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_330_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_349_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_349_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_349_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_349_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_349_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_349_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_368_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_368_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_368_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_368_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_368_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_368_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_381_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_381_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_381_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_381_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_381_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_393_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_393_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_393_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_393_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_393_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_405_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_405_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_405_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_405_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_405_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_431_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_431_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_431_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_431_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_431_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_443_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_443_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_443_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_443_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_443_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_455_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_455_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_455_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_455_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_455_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_467_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_467_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_467_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_467_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_467_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_47_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_47_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_47_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_47_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_47_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_47_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_712_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_712_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_712_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_712_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_712_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_712_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_922_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_922_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_922_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_922_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_922_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_922_word_offset_0 : std_logic_vector(10 downto 0);
    signal shl100_680 : std_logic_vector(63 downto 0);
    signal shl106_698 : std_logic_vector(63 downto 0);
    signal shl132_800 : std_logic_vector(63 downto 0);
    signal shl138_818 : std_logic_vector(63 downto 0);
    signal shl144_836 : std_logic_vector(63 downto 0);
    signal shl150_854 : std_logic_vector(63 downto 0);
    signal shl156_872 : std_logic_vector(63 downto 0);
    signal shl162_890 : std_logic_vector(63 downto 0);
    signal shl168_908 : std_logic_vector(63 downto 0);
    signal shl76_608 : std_logic_vector(63 downto 0);
    signal shl82_626 : std_logic_vector(63 downto 0);
    signal shl88_644 : std_logic_vector(63 downto 0);
    signal shl94_662 : std_logic_vector(63 downto 0);
    signal shl_590 : std_logic_vector(63 downto 0);
    signal shr123184x_xmask_514 : std_logic_vector(63 downto 0);
    signal shr188x_xmask_493 : std_logic_vector(63 downto 0);
    signal tmp11_233 : std_logic_vector(31 downto 0);
    signal tmp12_737 : std_logic_vector(31 downto 0);
    signal tmp13_742 : std_logic_vector(31 downto 0);
    signal tmp14_747 : std_logic_vector(31 downto 0);
    signal tmp15_751 : std_logic_vector(63 downto 0);
    signal tmp16_757 : std_logic_vector(63 downto 0);
    signal tmp17_763 : std_logic_vector(0 downto 0);
    signal tmp1_123 : std_logic_vector(31 downto 0);
    signal tmp230_223 : std_logic_vector(63 downto 0);
    signal tmp235_113 : std_logic_vector(63 downto 0);
    signal tmp3_195 : std_logic_vector(63 downto 0);
    signal tmp47_382 : std_logic_vector(31 downto 0);
    signal tmp48_394 : std_logic_vector(31 downto 0);
    signal tmp49_406 : std_logic_vector(31 downto 0);
    signal tmp53_432 : std_logic_vector(31 downto 0);
    signal tmp54_444 : std_logic_vector(31 downto 0);
    signal tmp56_456 : std_logic_vector(31 downto 0);
    signal tmp58_468 : std_logic_vector(31 downto 0);
    signal tmp5_532 : std_logic_vector(31 downto 0);
    signal tmp6_537 : std_logic_vector(31 downto 0);
    signal tmp7_541 : std_logic_vector(63 downto 0);
    signal tmp8_547 : std_logic_vector(63 downto 0);
    signal tmp9_553 : std_logic_vector(0 downto 0);
    signal tmp_92 : std_logic_vector(63 downto 0);
    signal type_cast_111_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_146_wire : std_logic_vector(31 downto 0);
    signal type_cast_153_wire : std_logic_vector(31 downto 0);
    signal type_cast_155_wire : std_logic_vector(31 downto 0);
    signal type_cast_170_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_185_wire : std_logic_vector(63 downto 0);
    signal type_cast_188_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_193_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_221_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_261_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_263_wire : std_logic_vector(63 downto 0);
    signal type_cast_267_wire : std_logic_vector(15 downto 0);
    signal type_cast_269_wire : std_logic_vector(15 downto 0);
    signal type_cast_290_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_296_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_309_wire : std_logic_vector(15 downto 0);
    signal type_cast_491_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_497_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_512_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_518_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_53_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_545_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_551_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_558_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_567_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_569_wire : std_logic_vector(63 downto 0);
    signal type_cast_588_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_606_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_624_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_642_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_660_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_678_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_696_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_718_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_755_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_761_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_768_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_76_wire : std_logic_vector(63 downto 0);
    signal type_cast_777_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_779_wire : std_logic_vector(63 downto 0);
    signal type_cast_798_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_79_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_816_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_834_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_83_wire : std_logic_vector(31 downto 0);
    signal type_cast_852_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_85_wire : std_logic_vector(31 downto 0);
    signal type_cast_870_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_888_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_906_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_90_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_928_wire_constant : std_logic_vector(63 downto 0);
    signal umax10_560 : std_logic_vector(63 downto 0);
    signal umax18_770 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_padding_311_word_address_0 <= "0";
    array_obj_ref_101_constant_part_of_offset <= "0000010";
    array_obj_ref_101_offset_scale_factor_0 <= "1000000";
    array_obj_ref_101_offset_scale_factor_1 <= "0000001";
    array_obj_ref_101_resized_base_address <= "0000000";
    array_obj_ref_204_constant_part_of_offset <= "0000010";
    array_obj_ref_204_offset_scale_factor_0 <= "1000000";
    array_obj_ref_204_offset_scale_factor_1 <= "0000001";
    array_obj_ref_204_resized_base_address <= "0000000";
    array_obj_ref_273_offset_scale_factor_0 <= "1";
    array_obj_ref_273_resized_base_address <= "0";
    array_obj_ref_575_constant_part_of_offset <= "00000000000000";
    array_obj_ref_575_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_575_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_575_resized_base_address <= "00000000000000";
    array_obj_ref_785_constant_part_of_offset <= "00000100001";
    array_obj_ref_785_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_785_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_785_resized_base_address <= "00000000000";
    iNsTr_13_119 <= "00000000000000000000000000000001";
    iNsTr_1_45 <= "00000000000000000000000000000001";
    iNsTr_21_229 <= "00000000000000000000000000000001";
    iNsTr_26_328 <= "00000000000000000000000000000010";
    iNsTr_29_347 <= "00000000000000000000000000000011";
    iNsTr_32_366 <= "00000000000000000000000000000100";
    iNsTr_34_378 <= "00000000000000000000000000000010";
    iNsTr_35_390 <= "00000000000000000000000000000011";
    iNsTr_36_402 <= "00000000000000000000000000000100";
    iNsTr_37_428 <= "00000000000000000000000000000010";
    iNsTr_38_440 <= "00000000000000000000000000000011";
    iNsTr_39_452 <= "00000000000000000000000000000100";
    iNsTr_40_464 <= "00000000000000000000000000000101";
    iNsTr_5_162 <= "00000000000000000000000000000001";
    ptr_deref_105_word_offset_0 <= "0000000";
    ptr_deref_122_word_offset_0 <= "0000000";
    ptr_deref_164_word_offset_0 <= "0000000";
    ptr_deref_215_word_offset_0 <= "0000000";
    ptr_deref_232_word_offset_0 <= "0000000";
    ptr_deref_277_word_offset_0 <= "0";
    ptr_deref_330_word_offset_0 <= "0000000";
    ptr_deref_349_word_offset_0 <= "0000000";
    ptr_deref_368_word_offset_0 <= "0000000";
    ptr_deref_381_word_offset_0 <= "0000000";
    ptr_deref_393_word_offset_0 <= "0000000";
    ptr_deref_405_word_offset_0 <= "0000000";
    ptr_deref_431_word_offset_0 <= "0000000";
    ptr_deref_443_word_offset_0 <= "0000000";
    ptr_deref_455_word_offset_0 <= "0000000";
    ptr_deref_467_word_offset_0 <= "0000000";
    ptr_deref_47_word_offset_0 <= "0000000";
    ptr_deref_712_word_offset_0 <= "00000000000000";
    ptr_deref_922_word_offset_0 <= "00000000000";
    type_cast_111_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_170_wire_constant <= "00000000000000000000000000000000";
    type_cast_188_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_193_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_221_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_261_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_290_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_296_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_491_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_497_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_512_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_518_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_53_wire_constant <= "00000000";
    type_cast_545_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_551_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_558_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_567_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_588_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_606_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_624_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_642_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_660_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_678_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_696_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_718_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_755_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_761_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_768_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_777_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_798_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_79_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_816_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_834_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_852_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_870_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_888_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_906_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_90_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_928_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_143: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_146_wire;
      req(0) <= phi_stmt_143_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_143",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_143_ack_0,
          idata => idata,
          odata => conv4x_xlcssa1_143,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_143
    phi_stmt_150: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_153_wire & type_cast_155_wire;
      req <= phi_stmt_150_req_0 & phi_stmt_150_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_150",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_150_ack_0,
          idata => idata,
          odata => conv4x_xlcssa_150,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_150
    phi_stmt_182: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_185_wire & type_cast_188_wire_constant;
      req <= phi_stmt_182_req_0 & phi_stmt_182_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_182",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_182_ack_0,
          idata => idata,
          odata => indvar228_182,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_182
    phi_stmt_257: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_261_wire_constant & type_cast_263_wire;
      req <= phi_stmt_257_req_0 & phi_stmt_257_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_257",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_257_ack_0,
          idata => idata,
          odata => indvar225_257,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_257
    phi_stmt_264: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_267_wire & type_cast_269_wire;
      req <= phi_stmt_264_req_0 & phi_stmt_264_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_264",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_264_ack_0,
          idata => idata,
          odata => conv30196_264,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_264
    phi_stmt_306: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_309_wire;
      req(0) <= phi_stmt_306_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_306",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_306_ack_0,
          idata => idata,
          odata => conv30x_xlcssa_306,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_306
    phi_stmt_563: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_567_wire_constant & type_cast_569_wire;
      req <= phi_stmt_563_req_0 & phi_stmt_563_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_563",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_563_ack_0,
          idata => idata,
          odata => indvar215_563,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_563
    phi_stmt_73: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_76_wire & type_cast_79_wire_constant;
      req <= phi_stmt_73_req_0 & phi_stmt_73_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_73",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_73_ack_0,
          idata => idata,
          odata => indvar233_73,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_73
    phi_stmt_773: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_777_wire_constant & type_cast_779_wire;
      req <= phi_stmt_773_req_0 & phi_stmt_773_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_773",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_773_ack_0,
          idata => idata,
          odata => indvar_773,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_773
    phi_stmt_80: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_83_wire & type_cast_85_wire;
      req <= phi_stmt_80_req_0 & phi_stmt_80_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_80",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_80_ack_0,
          idata => idata,
          odata => conv4207_80,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_80
    -- flow-through select operator MUX_559_inst
    umax10_560 <= tmp8_547 when (tmp9_553(0) /=  '0') else type_cast_558_wire_constant;
    -- flow-through select operator MUX_769_inst
    umax18_770 <= tmp16_757 when (tmp17_763(0) /=  '0') else type_cast_768_wire_constant;
    addr_of_102_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_102_final_reg_req_0;
      addr_of_102_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_102_final_reg_req_1;
      addr_of_102_final_reg_ack_1<= rack(0);
      addr_of_102_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_102_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_101_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_205_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_205_final_reg_req_0;
      addr_of_205_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_205_final_reg_req_1;
      addr_of_205_final_reg_ack_1<= rack(0);
      addr_of_205_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_205_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_204_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx19_206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_274_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_274_final_reg_req_0;
      addr_of_274_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_274_final_reg_req_1;
      addr_of_274_final_reg_ack_1<= rack(0);
      addr_of_274_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_274_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_273_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx33_275,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_576_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_576_final_reg_req_0;
      addr_of_576_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_576_final_reg_req_1;
      addr_of_576_final_reg_ack_1<= rack(0);
      addr_of_576_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_576_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_575_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx114_577,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_786_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_786_final_reg_req_0;
      addr_of_786_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_786_final_reg_req_1;
      addr_of_786_final_reg_ack_1<= rack(0);
      addr_of_786_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_786_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_785_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx176_787,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_134_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_134_inst_req_0;
      type_cast_134_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_134_inst_req_1;
      type_cast_134_inst_ack_1<= rack(0);
      type_cast_134_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_134_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_131,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_146_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_146_inst_req_0;
      type_cast_146_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_146_inst_req_1;
      type_cast_146_inst_ack_1<= rack(0);
      type_cast_146_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_146_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_146_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_153_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_153_inst_req_0;
      type_cast_153_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_153_inst_req_1;
      type_cast_153_inst_ack_1<= rack(0);
      type_cast_153_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_153_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4205_63,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_153_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_155_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_155_inst_req_0;
      type_cast_155_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_155_inst_req_1;
      type_cast_155_inst_ack_1<= rack(0);
      type_cast_155_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_155_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4x_xlcssa1_143,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_155_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_185_inst_req_0;
      type_cast_185_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_185_inst_req_1;
      type_cast_185_inst_ack_1<= rack(0);
      type_cast_185_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_185_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp230_223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_185_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_198_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_198_inst_req_0;
      type_cast_198_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_198_inst_req_1;
      type_cast_198_inst_ack_1<= rack(0);
      type_cast_198_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_198_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_195,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc22_199,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_212_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_212_inst_req_0;
      type_cast_212_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_212_inst_req_1;
      type_cast_212_inst_ack_1<= rack(0);
      type_cast_212_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_212_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_209,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_253_inst_req_0;
      type_cast_253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_253_inst_req_1;
      type_cast_253_inst_ack_1<= rack(0);
      type_cast_253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call29193_250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30194_254,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_263_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_263_inst_req_0;
      type_cast_263_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_263_inst_req_1;
      type_cast_263_inst_ack_1<= rack(0);
      type_cast_263_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_263_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext226_292,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_263_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_267_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_267_inst_req_0;
      type_cast_267_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_267_inst_req_1;
      type_cast_267_inst_ack_1<= rack(0);
      type_cast_267_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_267_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv30194_254,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_267_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_269_inst_req_0;
      type_cast_269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_269_inst_req_1;
      type_cast_269_inst_ack_1<= rack(0);
      type_cast_269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv30_286,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_269_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_285_inst_req_0;
      type_cast_285_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_285_inst_req_1;
      type_cast_285_inst_ack_1<= rack(0);
      type_cast_285_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_285_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call29_282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_286,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_309_inst_req_0;
      type_cast_309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_309_inst_req_1;
      type_cast_309_inst_ack_1<= rack(0);
      type_cast_309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv30_286,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_309_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_319_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_319_inst_req_0;
      type_cast_319_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_319_inst_req_1;
      type_cast_319_inst_ack_1<= rack(0);
      type_cast_319_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_319_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call40_316,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv41_320,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_338_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_338_inst_req_0;
      type_cast_338_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_338_inst_req_1;
      type_cast_338_inst_ack_1<= rack(0);
      type_cast_338_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_338_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call42_335,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv43_339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_357_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_357_inst_req_0;
      type_cast_357_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_357_inst_req_1;
      type_cast_357_inst_ack_1<= rack(0);
      type_cast_357_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_357_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call44_354,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv45_358,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_38_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_38_inst_req_0;
      type_cast_38_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_38_inst_req_1;
      type_cast_38_inst_ack_1<= rack(0);
      type_cast_38_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_38_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_39,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_419_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_419_inst_req_0;
      type_cast_419_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_419_inst_req_1;
      type_cast_419_inst_ack_1<= rack(0);
      type_cast_419_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_419_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul50_416,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_420,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_486_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_486_inst_req_0;
      type_cast_486_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_486_inst_req_1;
      type_cast_486_inst_ack_1<= rack(0);
      type_cast_486_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_486_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul59_483,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_487,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_540_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_540_inst_req_0;
      type_cast_540_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_540_inst_req_1;
      type_cast_540_inst_ack_1<= rack(0);
      type_cast_540_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_540_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp6_537,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp7_541,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_569_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_569_inst_req_0;
      type_cast_569_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_569_inst_req_1;
      type_cast_569_inst_ack_1<= rack(0);
      type_cast_569_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_569_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext216_720,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_569_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_583_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_583_inst_req_0;
      type_cast_583_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_583_inst_req_1;
      type_cast_583_inst_ack_1<= rack(0);
      type_cast_583_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_583_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call69_580,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_584,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_596_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_596_inst_req_0;
      type_cast_596_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_596_inst_req_1;
      type_cast_596_inst_ack_1<= rack(0);
      type_cast_596_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_596_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call72_593,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_597,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_614_inst_req_0;
      type_cast_614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_614_inst_req_1;
      type_cast_614_inst_ack_1<= rack(0);
      type_cast_614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call77_611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_62_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_62_inst_req_0;
      type_cast_62_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_62_inst_req_1;
      type_cast_62_inst_ack_1<= rack(0);
      type_cast_62_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_62_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3204_59,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4205_63,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_632_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_632_inst_req_0;
      type_cast_632_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_632_inst_req_1;
      type_cast_632_inst_ack_1<= rack(0);
      type_cast_632_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_632_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call83_629,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_633,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_650_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_650_inst_req_0;
      type_cast_650_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_650_inst_req_1;
      type_cast_650_inst_ack_1<= rack(0);
      type_cast_650_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_650_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_647,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_651,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_668_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_668_inst_req_0;
      type_cast_668_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_668_inst_req_1;
      type_cast_668_inst_ack_1<= rack(0);
      type_cast_668_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_668_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call95_665,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv97_669,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_686_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_686_inst_req_0;
      type_cast_686_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_686_inst_req_1;
      type_cast_686_inst_ack_1<= rack(0);
      type_cast_686_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_686_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_683,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv103_687,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_704_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_704_inst_req_0;
      type_cast_704_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_704_inst_req_1;
      type_cast_704_inst_ack_1<= rack(0);
      type_cast_704_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_704_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call107_701,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv109_705,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_750_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_750_inst_req_0;
      type_cast_750_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_750_inst_req_1;
      type_cast_750_inst_ack_1<= rack(0);
      type_cast_750_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_750_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp14_747,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_751,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_76_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_76_inst_req_0;
      type_cast_76_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_76_inst_req_1;
      type_cast_76_inst_ack_1<= rack(0);
      type_cast_76_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_76_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp235_113,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_76_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_779_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_779_inst_req_0;
      type_cast_779_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_779_inst_req_1;
      type_cast_779_inst_ack_1<= rack(0);
      type_cast_779_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_779_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_930,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_779_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_793_inst_req_0;
      type_cast_793_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_793_inst_req_1;
      type_cast_793_inst_ack_1<= rack(0);
      type_cast_793_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_793_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_790,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_794,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_806_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_806_inst_req_0;
      type_cast_806_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_806_inst_req_1;
      type_cast_806_inst_ack_1<= rack(0);
      type_cast_806_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_806_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_803,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv135_807,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_824_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_824_inst_req_0;
      type_cast_824_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_824_inst_req_1;
      type_cast_824_inst_ack_1<= rack(0);
      type_cast_824_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_824_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call139_821,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv141_825,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_83_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_83_inst_req_0;
      type_cast_83_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_83_inst_req_1;
      type_cast_83_inst_ack_1<= rack(0);
      type_cast_83_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_83_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_83_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_842_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_842_inst_req_0;
      type_cast_842_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_842_inst_req_1;
      type_cast_842_inst_ack_1<= rack(0);
      type_cast_842_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_842_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call145_839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_843,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_85_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_85_inst_req_0;
      type_cast_85_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_85_inst_req_1;
      type_cast_85_inst_ack_1<= rack(0);
      type_cast_85_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_85_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4205_63,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_85_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_860_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_860_inst_req_0;
      type_cast_860_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_860_inst_req_1;
      type_cast_860_inst_ack_1<= rack(0);
      type_cast_860_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_860_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call151_857,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_861,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_878_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_878_inst_req_0;
      type_cast_878_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_878_inst_req_1;
      type_cast_878_inst_ack_1<= rack(0);
      type_cast_878_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_878_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call157_875,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv159_879,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_896_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_896_inst_req_0;
      type_cast_896_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_896_inst_req_1;
      type_cast_896_inst_ack_1<= rack(0);
      type_cast_896_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_896_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call163_893,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_897,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_914_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_914_inst_req_0;
      type_cast_914_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_914_inst_req_1;
      type_cast_914_inst_ack_1<= rack(0);
      type_cast_914_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_914_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call169_911,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv171_915,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_947_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_947_inst_req_0;
      type_cast_947_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_947_inst_req_1;
      type_cast_947_inst_ack_1<= rack(0);
      type_cast_947_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_947_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul50_416,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ret_val_x_x_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_95_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_95_inst_req_0;
      type_cast_95_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_95_inst_req_1;
      type_cast_95_inst_ack_1<= rack(0);
      type_cast_95_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_95_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_92,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc_96,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_padding_311_gather_scatter
    process(conv30x_xlcssa_306) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv30x_xlcssa_306;
      ov(15 downto 0) := iv;
      STORE_padding_311_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_index_1_rename
    process(R_indvar233_100_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar233_100_resized;
      ov(6 downto 0) := iv;
      R_indvar233_100_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_index_1_resize
    process(indvar233_73) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar233_73;
      ov := iv(6 downto 0);
      R_indvar233_100_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_root_address_inst
    process(array_obj_ref_101_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_101_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_101_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_204_index_1_rename
    process(R_indvar228_203_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar228_203_resized;
      ov(6 downto 0) := iv;
      R_indvar228_203_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_204_index_1_resize
    process(indvar228_182) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar228_182;
      ov := iv(6 downto 0);
      R_indvar228_203_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_204_root_address_inst
    process(array_obj_ref_204_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_204_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_204_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_273_index_0_rename
    process(R_indvar225_272_resized) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar225_272_resized;
      ov(0 downto 0) := iv;
      R_indvar225_272_scaled <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_273_index_0_resize
    process(indvar225_257) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar225_257;
      ov := iv(0 downto 0);
      R_indvar225_272_resized <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_273_index_offset
    process(R_indvar225_272_scaled) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar225_272_scaled;
      ov(0 downto 0) := iv;
      array_obj_ref_273_final_offset <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_273_root_address_inst
    process(array_obj_ref_273_final_offset) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_273_final_offset;
      ov(0 downto 0) := iv;
      array_obj_ref_273_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_575_index_1_rename
    process(R_indvar215_574_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar215_574_resized;
      ov(13 downto 0) := iv;
      R_indvar215_574_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_575_index_1_resize
    process(indvar215_563) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar215_563;
      ov := iv(13 downto 0);
      R_indvar215_574_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_575_root_address_inst
    process(array_obj_ref_575_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_575_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_575_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_785_index_1_rename
    process(R_indvar_784_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_784_resized;
      ov(10 downto 0) := iv;
      R_indvar_784_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_785_index_1_resize
    process(indvar_773) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_773;
      ov := iv(10 downto 0);
      R_indvar_784_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_785_root_address_inst
    process(array_obj_ref_785_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_785_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_785_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_addr_0
    process(ptr_deref_105_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_105_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_105_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_base_resize
    process(arrayidx_103) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_103;
      ov := iv(6 downto 0);
      ptr_deref_105_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_gather_scatter
    process(conv4207_80) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv4207_80;
      ov(31 downto 0) := iv;
      ptr_deref_105_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_root_address_inst
    process(ptr_deref_105_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_105_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_105_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_addr_0
    process(ptr_deref_122_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_122_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_122_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_base_resize
    process(iNsTr_13_119) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_13_119;
      ov := iv(6 downto 0);
      ptr_deref_122_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_gather_scatter
    process(ptr_deref_122_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_122_data_0;
      ov(31 downto 0) := iv;
      tmp1_123 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_root_address_inst
    process(ptr_deref_122_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_122_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_122_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_164_addr_0
    process(ptr_deref_164_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_164_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_164_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_164_base_resize
    process(iNsTr_5_162) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_162;
      ov := iv(6 downto 0);
      ptr_deref_164_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_164_gather_scatter
    process(conv4x_xlcssa_150) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv4x_xlcssa_150;
      ov(31 downto 0) := iv;
      ptr_deref_164_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_164_root_address_inst
    process(ptr_deref_164_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_164_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_164_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_215_addr_0
    process(ptr_deref_215_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_215_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_215_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_215_base_resize
    process(arrayidx19_206) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx19_206;
      ov := iv(6 downto 0);
      ptr_deref_215_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_215_gather_scatter
    process(conv16_213) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv16_213;
      ov(31 downto 0) := iv;
      ptr_deref_215_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_215_root_address_inst
    process(ptr_deref_215_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_215_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_215_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_232_addr_0
    process(ptr_deref_232_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_232_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_232_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_232_base_resize
    process(iNsTr_21_229) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_21_229;
      ov := iv(6 downto 0);
      ptr_deref_232_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_232_gather_scatter
    process(ptr_deref_232_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_232_data_0;
      ov(31 downto 0) := iv;
      tmp11_233 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_232_root_address_inst
    process(ptr_deref_232_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_232_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_232_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_277_addr_0
    process(ptr_deref_277_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_277_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_277_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_277_base_resize
    process(arrayidx33_275) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx33_275;
      ov := iv(0 downto 0);
      ptr_deref_277_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_277_gather_scatter
    process(conv30196_264) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv30196_264;
      ov(15 downto 0) := iv;
      ptr_deref_277_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_277_root_address_inst
    process(ptr_deref_277_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_277_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_277_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_330_addr_0
    process(ptr_deref_330_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_330_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_330_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_330_base_resize
    process(iNsTr_26_328) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_26_328;
      ov := iv(6 downto 0);
      ptr_deref_330_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_330_gather_scatter
    process(conv41_320) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv41_320;
      ov(31 downto 0) := iv;
      ptr_deref_330_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_330_root_address_inst
    process(ptr_deref_330_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_330_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_330_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_349_addr_0
    process(ptr_deref_349_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_349_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_349_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_349_base_resize
    process(iNsTr_29_347) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_29_347;
      ov := iv(6 downto 0);
      ptr_deref_349_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_349_gather_scatter
    process(conv43_339) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv43_339;
      ov(31 downto 0) := iv;
      ptr_deref_349_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_349_root_address_inst
    process(ptr_deref_349_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_349_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_349_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_368_addr_0
    process(ptr_deref_368_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_368_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_368_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_368_base_resize
    process(iNsTr_32_366) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_32_366;
      ov := iv(6 downto 0);
      ptr_deref_368_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_368_gather_scatter
    process(conv45_358) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv45_358;
      ov(31 downto 0) := iv;
      ptr_deref_368_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_368_root_address_inst
    process(ptr_deref_368_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_368_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_368_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_addr_0
    process(ptr_deref_381_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_381_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_381_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_base_resize
    process(iNsTr_34_378) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_34_378;
      ov := iv(6 downto 0);
      ptr_deref_381_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_gather_scatter
    process(ptr_deref_381_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_381_data_0;
      ov(31 downto 0) := iv;
      tmp47_382 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_root_address_inst
    process(ptr_deref_381_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_381_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_381_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_393_addr_0
    process(ptr_deref_393_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_393_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_393_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_393_base_resize
    process(iNsTr_35_390) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_35_390;
      ov := iv(6 downto 0);
      ptr_deref_393_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_393_gather_scatter
    process(ptr_deref_393_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_393_data_0;
      ov(31 downto 0) := iv;
      tmp48_394 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_393_root_address_inst
    process(ptr_deref_393_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_393_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_393_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_405_addr_0
    process(ptr_deref_405_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_405_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_405_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_405_base_resize
    process(iNsTr_36_402) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_36_402;
      ov := iv(6 downto 0);
      ptr_deref_405_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_405_gather_scatter
    process(ptr_deref_405_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_405_data_0;
      ov(31 downto 0) := iv;
      tmp49_406 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_405_root_address_inst
    process(ptr_deref_405_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_405_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_405_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_431_addr_0
    process(ptr_deref_431_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_431_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_431_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_431_base_resize
    process(iNsTr_37_428) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_37_428;
      ov := iv(6 downto 0);
      ptr_deref_431_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_431_gather_scatter
    process(ptr_deref_431_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_431_data_0;
      ov(31 downto 0) := iv;
      tmp53_432 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_431_root_address_inst
    process(ptr_deref_431_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_431_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_431_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_443_addr_0
    process(ptr_deref_443_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_443_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_443_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_443_base_resize
    process(iNsTr_38_440) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_38_440;
      ov := iv(6 downto 0);
      ptr_deref_443_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_443_gather_scatter
    process(ptr_deref_443_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_443_data_0;
      ov(31 downto 0) := iv;
      tmp54_444 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_443_root_address_inst
    process(ptr_deref_443_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_443_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_443_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_455_addr_0
    process(ptr_deref_455_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_455_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_455_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_455_base_resize
    process(iNsTr_39_452) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_39_452;
      ov := iv(6 downto 0);
      ptr_deref_455_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_455_gather_scatter
    process(ptr_deref_455_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_455_data_0;
      ov(31 downto 0) := iv;
      tmp56_456 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_455_root_address_inst
    process(ptr_deref_455_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_455_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_455_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_467_addr_0
    process(ptr_deref_467_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_467_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_467_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_467_base_resize
    process(iNsTr_40_464) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_40_464;
      ov := iv(6 downto 0);
      ptr_deref_467_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_467_gather_scatter
    process(ptr_deref_467_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_467_data_0;
      ov(31 downto 0) := iv;
      tmp58_468 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_467_root_address_inst
    process(ptr_deref_467_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_467_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_467_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_addr_0
    process(ptr_deref_47_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_47_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_47_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_base_resize
    process(iNsTr_1_45) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_45;
      ov := iv(6 downto 0);
      ptr_deref_47_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_gather_scatter
    process(conv_39) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_39;
      ov(31 downto 0) := iv;
      ptr_deref_47_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_root_address_inst
    process(ptr_deref_47_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_47_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_47_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_712_addr_0
    process(ptr_deref_712_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_712_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_712_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_712_base_resize
    process(arrayidx114_577) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx114_577;
      ov := iv(13 downto 0);
      ptr_deref_712_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_712_gather_scatter
    process(add110_710) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add110_710;
      ov(63 downto 0) := iv;
      ptr_deref_712_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_712_root_address_inst
    process(ptr_deref_712_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_712_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_712_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_922_addr_0
    process(ptr_deref_922_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_922_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_922_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_922_base_resize
    process(arrayidx176_787) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx176_787;
      ov := iv(10 downto 0);
      ptr_deref_922_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_922_gather_scatter
    process(add172_920) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add172_920;
      ov(63 downto 0) := iv;
      ptr_deref_922_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_922_root_address_inst
    process(ptr_deref_922_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_922_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_922_root_address <= ov(10 downto 0);
      --
    end process;
    if_stmt_136_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_128;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_136_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_136_branch_req_0,
          ack0 => if_stmt_136_branch_ack_0,
          ack1 => if_stmt_136_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_173_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp12199_172;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_173_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_173_branch_req_0,
          ack0 => if_stmt_173_branch_ack_0,
          ack1 => if_stmt_173_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_239_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp12_238;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_239_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_239_branch_req_0,
          ack0 => if_stmt_239_branch_ack_0,
          ack1 => if_stmt_239_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_299_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_298;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_299_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_299_branch_req_0,
          ack0 => if_stmt_299_branch_ack_0,
          ack1 => if_stmt_299_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_500_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp65189_499;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_500_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_500_branch_req_0,
          ack0 => if_stmt_500_branch_ack_0,
          ack1 => if_stmt_500_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_521_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp124185_520;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_521_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_521_branch_req_0,
          ack0 => if_stmt_521_branch_ack_0,
          ack1 => if_stmt_521_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_64_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp203_56;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_64_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_64_branch_req_0,
          ack0 => if_stmt_64_branch_ack_0,
          ack1 => if_stmt_64_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_726_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond11_725;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_726_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_726_branch_req_0,
          ack0 => if_stmt_726_branch_ack_0,
          ack1 => if_stmt_726_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_936_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond19_935;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_936_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_936_branch_req_0,
          ack0 => if_stmt_936_branch_ack_0,
          ack1 => if_stmt_936_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_112_inst
    process(indvar233_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar233_73, type_cast_111_wire_constant, tmp_var);
      tmp235_113 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_194_inst
    process(indvar228_182) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar228_182, type_cast_193_wire_constant, tmp_var);
      tmp3_195 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_222_inst
    process(indvar228_182) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar228_182, type_cast_221_wire_constant, tmp_var);
      tmp230_223 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_291_inst
    process(indvar225_257) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar225_257, type_cast_290_wire_constant, tmp_var);
      indvarx_xnext226_292 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_719_inst
    process(indvar215_563) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar215_563, type_cast_718_wire_constant, tmp_var);
      indvarx_xnext216_720 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_91_inst
    process(indvar233_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar233_73, type_cast_90_wire_constant, tmp_var);
      tmp_92 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_929_inst
    process(indvar_773) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_773, type_cast_928_wire_constant, tmp_var);
      indvarx_xnext_930 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_492_inst
    process(conv51_420) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv51_420, type_cast_491_wire_constant, tmp_var);
      shr188x_xmask_493 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_513_inst
    process(conv60_487) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv60_487, type_cast_512_wire_constant, tmp_var);
      shr123184x_xmask_514 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_171_inst
    process(conv4x_xlcssa_150) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv4x_xlcssa_150, type_cast_170_wire_constant, tmp_var);
      cmp12199_172 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_297_inst
    process(indvarx_xnext226_292) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext226_292, type_cast_296_wire_constant, tmp_var);
      exitcond_298 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_498_inst
    process(shr188x_xmask_493) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr188x_xmask_493, type_cast_497_wire_constant, tmp_var);
      cmp65189_499 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_519_inst
    process(shr123184x_xmask_514) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr123184x_xmask_514, type_cast_518_wire_constant, tmp_var);
      cmp124185_520 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_724_inst
    process(indvarx_xnext216_720, umax10_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext216_720, umax10_560, tmp_var);
      exitcond11_725 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_934_inst
    process(indvarx_xnext_930, umax18_770) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_930, umax18_770, tmp_var);
      exitcond19_935 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_54_inst
    process(call_35) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(call_35, type_cast_53_wire_constant, tmp_var);
      cmp203_56 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_546_inst
    process(tmp7_541) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp7_541, type_cast_545_wire_constant, tmp_var);
      tmp8_547 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_756_inst
    process(tmp15_751) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp15_751, type_cast_755_wire_constant, tmp_var);
      tmp16_757 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_410_inst
    process(tmp48_394, tmp47_382) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp48_394, tmp47_382, tmp_var);
      mul_411 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_415_inst
    process(mul_411, tmp49_406) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_411, tmp49_406, tmp_var);
      mul50_416 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_472_inst
    process(tmp54_444, tmp53_432) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_444, tmp53_432, tmp_var);
      mul55_473 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_477_inst
    process(mul55_473, tmp56_456) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul55_473, tmp56_456, tmp_var);
      mul57_478 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_482_inst
    process(mul57_478, tmp58_468) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul57_478, tmp58_468, tmp_var);
      mul59_483 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_531_inst
    process(tmp48_394, tmp47_382) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp48_394, tmp47_382, tmp_var);
      tmp5_532 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_536_inst
    process(tmp5_532, tmp49_406) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp5_532, tmp49_406, tmp_var);
      tmp6_537 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_736_inst
    process(tmp54_444, tmp53_432) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_444, tmp53_432, tmp_var);
      tmp12_737 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_741_inst
    process(tmp12_737, tmp56_456) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_737, tmp56_456, tmp_var);
      tmp13_742 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_746_inst
    process(tmp13_742, tmp58_468) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp13_742, tmp58_468, tmp_var);
      tmp14_747 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_601_inst
    process(shl_590, conv74_597) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_590, conv74_597, tmp_var);
      add_602 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_619_inst
    process(shl76_608, conv79_615) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl76_608, conv79_615, tmp_var);
      add80_620 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_637_inst
    process(shl82_626, conv85_633) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl82_626, conv85_633, tmp_var);
      add86_638 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_655_inst
    process(shl88_644, conv91_651) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl88_644, conv91_651, tmp_var);
      add92_656 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_673_inst
    process(shl94_662, conv97_669) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl94_662, conv97_669, tmp_var);
      add98_674 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_691_inst
    process(shl100_680, conv103_687) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl100_680, conv103_687, tmp_var);
      add104_692 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_709_inst
    process(shl106_698, conv109_705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl106_698, conv109_705, tmp_var);
      add110_710 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_811_inst
    process(shl132_800, conv135_807) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_800, conv135_807, tmp_var);
      add136_812 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_829_inst
    process(shl138_818, conv141_825) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl138_818, conv141_825, tmp_var);
      add142_830 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_847_inst
    process(shl144_836, conv147_843) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl144_836, conv147_843, tmp_var);
      add148_848 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_865_inst
    process(shl150_854, conv153_861) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl150_854, conv153_861, tmp_var);
      add154_866 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_883_inst
    process(shl156_872, conv159_879) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl156_872, conv159_879, tmp_var);
      add160_884 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_901_inst
    process(shl162_890, conv165_897) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl162_890, conv165_897, tmp_var);
      add166_902 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_919_inst
    process(shl168_908, conv171_915) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl168_908, conv171_915, tmp_var);
      add172_920 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_589_inst
    process(conv70_584) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv70_584, type_cast_588_wire_constant, tmp_var);
      shl_590 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_607_inst
    process(add_602) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_602, type_cast_606_wire_constant, tmp_var);
      shl76_608 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_625_inst
    process(add80_620) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add80_620, type_cast_624_wire_constant, tmp_var);
      shl82_626 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_643_inst
    process(add86_638) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add86_638, type_cast_642_wire_constant, tmp_var);
      shl88_644 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_661_inst
    process(add92_656) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add92_656, type_cast_660_wire_constant, tmp_var);
      shl94_662 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_679_inst
    process(add98_674) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add98_674, type_cast_678_wire_constant, tmp_var);
      shl100_680 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_697_inst
    process(add104_692) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add104_692, type_cast_696_wire_constant, tmp_var);
      shl106_698 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_799_inst
    process(conv130_794) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv130_794, type_cast_798_wire_constant, tmp_var);
      shl132_800 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_817_inst
    process(add136_812) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add136_812, type_cast_816_wire_constant, tmp_var);
      shl138_818 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_835_inst
    process(add142_830) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add142_830, type_cast_834_wire_constant, tmp_var);
      shl144_836 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_853_inst
    process(add148_848) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add148_848, type_cast_852_wire_constant, tmp_var);
      shl150_854 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_871_inst
    process(add154_866) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add154_866, type_cast_870_wire_constant, tmp_var);
      shl156_872 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_889_inst
    process(add160_884) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add160_884, type_cast_888_wire_constant, tmp_var);
      shl162_890 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_907_inst
    process(add166_902) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add166_902, type_cast_906_wire_constant, tmp_var);
      shl168_908 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_552_inst
    process(tmp8_547) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp8_547, type_cast_551_wire_constant, tmp_var);
      tmp9_553 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_762_inst
    process(tmp16_757) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp16_757, type_cast_761_wire_constant, tmp_var);
      tmp17_763 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_127_inst
    process(inc_96, tmp1_123) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(inc_96, tmp1_123, tmp_var);
      cmp_128 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_237_inst
    process(inc22_199, tmp11_233) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(inc22_199, tmp11_233, tmp_var);
      cmp12_238 <= tmp_var; --
    end process;
    -- shared split operator group (60) : array_obj_ref_101_index_offset 
    ApIntAdd_group_60: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar233_100_scaled;
      array_obj_ref_101_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_101_index_offset_req_0;
      array_obj_ref_101_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_101_index_offset_req_1;
      array_obj_ref_101_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_60_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_60_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_60",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000010",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : array_obj_ref_204_index_offset 
    ApIntAdd_group_61: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar228_203_scaled;
      array_obj_ref_204_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_204_index_offset_req_0;
      array_obj_ref_204_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_204_index_offset_req_1;
      array_obj_ref_204_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_61_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_61_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_61",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000010",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : array_obj_ref_575_index_offset 
    ApIntAdd_group_62: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar215_574_scaled;
      array_obj_ref_575_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_575_index_offset_req_0;
      array_obj_ref_575_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_575_index_offset_req_1;
      array_obj_ref_575_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_62_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_62_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_62",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : array_obj_ref_785_index_offset 
    ApIntAdd_group_63: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_784_scaled;
      array_obj_ref_785_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_785_index_offset_req_0;
      array_obj_ref_785_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_785_index_offset_req_1;
      array_obj_ref_785_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_63_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_63_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_63",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100001",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared load operator group (0) : ptr_deref_122_load_0 ptr_deref_381_load_0 ptr_deref_393_load_0 ptr_deref_405_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_122_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_381_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_393_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_405_load_0_req_0;
      ptr_deref_122_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_381_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_393_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_405_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_122_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_381_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_393_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_405_load_0_req_1;
      ptr_deref_122_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_381_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_393_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_405_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_122_word_address_0 & ptr_deref_381_word_address_0 & ptr_deref_393_word_address_0 & ptr_deref_405_word_address_0;
      ptr_deref_122_data_0 <= data_out(127 downto 96);
      ptr_deref_381_data_0 <= data_out(95 downto 64);
      ptr_deref_393_data_0 <= data_out(63 downto 32);
      ptr_deref_405_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_232_load_0 ptr_deref_431_load_0 ptr_deref_443_load_0 ptr_deref_455_load_0 ptr_deref_467_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(34 downto 0);
      signal data_out: std_logic_vector(159 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant inBUFs : IntegerArray(4 downto 0) := (4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2);
      -- 
    begin -- 
      reqL_unguarded(4) <= ptr_deref_232_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_431_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_443_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_455_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_467_load_0_req_0;
      ptr_deref_232_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_431_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_443_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_455_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_467_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= ptr_deref_232_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_431_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_443_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_455_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_467_load_0_req_1;
      ptr_deref_232_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_431_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_443_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_455_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_467_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 5, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_232_word_address_0 & ptr_deref_431_word_address_0 & ptr_deref_443_word_address_0 & ptr_deref_455_word_address_0 & ptr_deref_467_word_address_0;
      ptr_deref_232_data_0 <= data_out(159 downto 128);
      ptr_deref_431_data_0 <= data_out(127 downto 96);
      ptr_deref_443_data_0 <= data_out(95 downto 64);
      ptr_deref_455_data_0 <= data_out(63 downto 32);
      ptr_deref_467_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 5,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 5,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared store operator group (0) : STORE_padding_311_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_padding_311_store_0_req_0;
      STORE_padding_311_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_padding_311_store_0_req_1;
      STORE_padding_311_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_padding_311_word_address_0;
      data_in <= STORE_padding_311_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(0 downto 0),
          mdata => memory_space_6_sr_data(15 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_105_store_0 ptr_deref_47_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_105_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_47_store_0_req_0;
      ptr_deref_105_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_47_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_105_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_47_store_0_req_1;
      ptr_deref_105_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_47_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_105_word_address_0 & ptr_deref_47_word_address_0;
      data_in <= ptr_deref_105_data_0 & ptr_deref_47_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(6 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_164_store_0 ptr_deref_215_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_164_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_215_store_0_req_0;
      ptr_deref_164_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_215_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_164_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_215_store_0_req_1;
      ptr_deref_164_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_215_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup2_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_164_word_address_0 & ptr_deref_215_word_address_0;
      data_in <= ptr_deref_164_data_0 & ptr_deref_215_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(6 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_277_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_277_store_0_req_0;
      ptr_deref_277_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_277_store_0_req_1;
      ptr_deref_277_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_277_word_address_0;
      data_in <= ptr_deref_277_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(15 downto 0),
          mtag => memory_space_7_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_330_store_0 ptr_deref_349_store_0 ptr_deref_368_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_330_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_349_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_368_store_0_req_0;
      ptr_deref_330_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_349_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_368_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_330_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_349_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_368_store_0_req_1;
      ptr_deref_330_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_349_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_368_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup4_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_330_word_address_0 & ptr_deref_349_word_address_0 & ptr_deref_368_word_address_0;
      data_in <= ptr_deref_330_data_0 & ptr_deref_349_data_0 & ptr_deref_368_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(6 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_712_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_712_store_0_req_0;
      ptr_deref_712_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_712_store_0_req_1;
      ptr_deref_712_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_712_word_address_0;
      data_in <= ptr_deref_712_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_922_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_922_store_0_req_0;
      ptr_deref_922_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_922_store_0_req_1;
      ptr_deref_922_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_922_word_address_0;
      data_in <= ptr_deref_922_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(10 downto 0),
          mdata => memory_space_4_sr_data(63 downto 0),
          mtag => memory_space_4_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared inport operator group (0) : RPIPE_ConvTranspose_input_pipe_58_inst RPIPE_ConvTranspose_input_pipe_34_inst RPIPE_ConvTranspose_input_pipe_130_inst RPIPE_ConvTranspose_input_pipe_353_inst RPIPE_ConvTranspose_input_pipe_315_inst RPIPE_ConvTranspose_input_pipe_281_inst RPIPE_ConvTranspose_input_pipe_892_inst RPIPE_ConvTranspose_input_pipe_249_inst RPIPE_ConvTranspose_input_pipe_334_inst RPIPE_ConvTranspose_input_pipe_910_inst RPIPE_ConvTranspose_input_pipe_208_inst RPIPE_ConvTranspose_input_pipe_579_inst RPIPE_ConvTranspose_input_pipe_592_inst RPIPE_ConvTranspose_input_pipe_874_inst RPIPE_ConvTranspose_input_pipe_610_inst RPIPE_ConvTranspose_input_pipe_856_inst RPIPE_ConvTranspose_input_pipe_628_inst RPIPE_ConvTranspose_input_pipe_838_inst RPIPE_ConvTranspose_input_pipe_646_inst RPIPE_ConvTranspose_input_pipe_820_inst RPIPE_ConvTranspose_input_pipe_664_inst RPIPE_ConvTranspose_input_pipe_802_inst RPIPE_ConvTranspose_input_pipe_682_inst RPIPE_ConvTranspose_input_pipe_789_inst RPIPE_ConvTranspose_input_pipe_700_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(199 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 24 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 24 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 24 downto 0);
      signal guard_vector : std_logic_vector( 24 downto 0);
      constant outBUFs : IntegerArray(24 downto 0) := (24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(24 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false);
      constant guardBuffering: IntegerArray(24 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2);
      -- 
    begin -- 
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_58_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_130_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_353_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_315_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_281_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_892_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_249_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_334_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_910_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_208_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_579_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_592_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_874_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_610_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_856_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_628_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_838_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_646_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_820_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_664_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_802_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_682_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_789_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_700_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_58_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_130_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_353_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_315_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_281_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_892_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_249_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_334_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_910_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_208_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_579_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_592_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_874_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_610_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_856_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_628_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_838_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_646_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_820_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_664_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_802_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_682_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_789_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_700_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_58_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_130_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_353_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_315_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_281_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_892_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_249_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_334_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_910_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_208_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_579_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_592_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_874_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_610_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_856_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_628_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_838_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_646_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_820_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_664_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_802_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_682_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_789_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_700_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_58_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_130_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_353_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_315_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_281_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_892_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_249_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_334_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_910_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_208_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_579_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_592_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_874_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_610_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_856_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_628_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_838_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_646_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_820_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_664_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_802_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_682_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_789_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_700_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      call3204_59 <= data_out(199 downto 192);
      call_35 <= data_out(191 downto 184);
      call3_131 <= data_out(183 downto 176);
      call44_354 <= data_out(175 downto 168);
      call40_316 <= data_out(167 downto 160);
      call29_282 <= data_out(159 downto 152);
      call163_893 <= data_out(151 downto 144);
      call29193_250 <= data_out(143 downto 136);
      call42_335 <= data_out(135 downto 128);
      call169_911 <= data_out(127 downto 120);
      call15_209 <= data_out(119 downto 112);
      call69_580 <= data_out(111 downto 104);
      call72_593 <= data_out(103 downto 96);
      call157_875 <= data_out(95 downto 88);
      call77_611 <= data_out(87 downto 80);
      call151_857 <= data_out(79 downto 72);
      call83_629 <= data_out(71 downto 64);
      call145_839 <= data_out(63 downto 56);
      call89_647 <= data_out(55 downto 48);
      call139_821 <= data_out(47 downto 40);
      call95_665 <= data_out(39 downto 32);
      call133_803 <= data_out(31 downto 24);
      call101_683 <= data_out(23 downto 16);
      call129_790 <= data_out(15 downto 8);
      call107_701 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_0_gI", nreqs => 25, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_0", data_width => 8,  num_reqs => 25,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(159 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(159 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(99 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(159 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(9 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(3 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(3 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(55 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(255 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(75 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(3 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(79 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_data : in   std_logic_vector(15 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal testConfigure_out_args   : std_logic_vector(15 downto 0);
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_data: std_logic_vector(15 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_data => testConfigure_return_data(15 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(3 downto 3),
      memory_space_0_lr_ack => memory_space_0_lr_ack(3 downto 3),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 21),
      memory_space_0_lr_tag => memory_space_0_lr_tag(83 downto 63),
      memory_space_0_lc_req => memory_space_0_lc_req(3 downto 3),
      memory_space_0_lc_ack => memory_space_0_lc_ack(3 downto 3),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 96),
      memory_space_0_lc_tag => memory_space_0_lc_tag(11 downto 9),
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 21),
      memory_space_1_lr_tag => memory_space_1_lr_tag(83 downto 63),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 96),
      memory_space_1_lc_tag => memory_space_1_lc_tag(11 downto 9),
      memory_space_2_lr_req => memory_space_2_lr_req(3 downto 3),
      memory_space_2_lr_ack => memory_space_2_lr_ack(3 downto 3),
      memory_space_2_lr_addr => memory_space_2_lr_addr(27 downto 21),
      memory_space_2_lr_tag => memory_space_2_lr_tag(79 downto 60),
      memory_space_2_lc_req => memory_space_2_lc_req(3 downto 3),
      memory_space_2_lc_ack => memory_space_2_lc_ack(3 downto 3),
      memory_space_2_lc_data => memory_space_2_lc_data(127 downto 96),
      memory_space_2_lc_tag => memory_space_2_lc_tag(7 downto 6),
      memory_space_3_lr_req => memory_space_3_lr_req(3 downto 3),
      memory_space_3_lr_ack => memory_space_3_lr_ack(3 downto 3),
      memory_space_3_lr_addr => memory_space_3_lr_addr(55 downto 42),
      memory_space_3_lr_tag => memory_space_3_lr_tag(75 downto 57),
      memory_space_3_lc_req => memory_space_3_lc_req(3 downto 3),
      memory_space_3_lc_ack => memory_space_3_lc_ack(3 downto 3),
      memory_space_3_lc_data => memory_space_3_lc_data(255 downto 192),
      memory_space_3_lc_tag => memory_space_3_lc_tag(3 downto 3),
      memory_space_6_lr_req => memory_space_6_lr_req(3 downto 3),
      memory_space_6_lr_ack => memory_space_6_lr_ack(3 downto 3),
      memory_space_6_lr_addr => memory_space_6_lr_addr(3 downto 3),
      memory_space_6_lr_tag => memory_space_6_lr_tag(75 downto 57),
      memory_space_6_lc_req => memory_space_6_lc_req(3 downto 3),
      memory_space_6_lc_ack => memory_space_6_lc_ack(3 downto 3),
      memory_space_6_lc_data => memory_space_6_lc_data(63 downto 48),
      memory_space_6_lc_tag => memory_space_6_lc_tag(3 downto 3),
      memory_space_7_lr_req => memory_space_7_lr_req(3 downto 3),
      memory_space_7_lr_ack => memory_space_7_lr_ack(3 downto 3),
      memory_space_7_lr_addr => memory_space_7_lr_addr(3 downto 3),
      memory_space_7_lr_tag => memory_space_7_lr_tag(79 downto 60),
      memory_space_7_lc_req => memory_space_7_lc_req(3 downto 3),
      memory_space_7_lc_ack => memory_space_7_lc_ack(3 downto 3),
      memory_space_7_lc_data => memory_space_7_lc_data(63 downto 48),
      memory_space_7_lc_tag => memory_space_7_lc_tag(7 downto 6),
      memory_space_5_sr_req => memory_space_5_sr_req(3 downto 3),
      memory_space_5_sr_ack => memory_space_5_sr_ack(3 downto 3),
      memory_space_5_sr_addr => memory_space_5_sr_addr(55 downto 42),
      memory_space_5_sr_data => memory_space_5_sr_data(255 downto 192),
      memory_space_5_sr_tag => memory_space_5_sr_tag(75 downto 57),
      memory_space_5_sc_req => memory_space_5_sc_req(3 downto 3),
      memory_space_5_sc_ack => memory_space_5_sc_ack(3 downto 3),
      memory_space_5_sc_tag => memory_space_5_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(2 downto 2),
      memory_space_0_lr_ack => memory_space_0_lr_ack(2 downto 2),
      memory_space_0_lr_addr => memory_space_0_lr_addr(20 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(62 downto 42),
      memory_space_0_lc_req => memory_space_0_lc_req(2 downto 2),
      memory_space_0_lc_ack => memory_space_0_lc_ack(2 downto 2),
      memory_space_0_lc_data => memory_space_0_lc_data(95 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(8 downto 6),
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(20 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(62 downto 42),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(95 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(8 downto 6),
      memory_space_2_lr_req => memory_space_2_lr_req(2 downto 2),
      memory_space_2_lr_ack => memory_space_2_lr_ack(2 downto 2),
      memory_space_2_lr_addr => memory_space_2_lr_addr(20 downto 14),
      memory_space_2_lr_tag => memory_space_2_lr_tag(59 downto 40),
      memory_space_2_lc_req => memory_space_2_lc_req(2 downto 2),
      memory_space_2_lc_ack => memory_space_2_lc_ack(2 downto 2),
      memory_space_2_lc_data => memory_space_2_lc_data(95 downto 64),
      memory_space_2_lc_tag => memory_space_2_lc_tag(5 downto 4),
      memory_space_3_lr_req => memory_space_3_lr_req(2 downto 2),
      memory_space_3_lr_ack => memory_space_3_lr_ack(2 downto 2),
      memory_space_3_lr_addr => memory_space_3_lr_addr(41 downto 28),
      memory_space_3_lr_tag => memory_space_3_lr_tag(56 downto 38),
      memory_space_3_lc_req => memory_space_3_lc_req(2 downto 2),
      memory_space_3_lc_ack => memory_space_3_lc_ack(2 downto 2),
      memory_space_3_lc_data => memory_space_3_lc_data(191 downto 128),
      memory_space_3_lc_tag => memory_space_3_lc_tag(2 downto 2),
      memory_space_6_lr_req => memory_space_6_lr_req(2 downto 2),
      memory_space_6_lr_ack => memory_space_6_lr_ack(2 downto 2),
      memory_space_6_lr_addr => memory_space_6_lr_addr(2 downto 2),
      memory_space_6_lr_tag => memory_space_6_lr_tag(56 downto 38),
      memory_space_6_lc_req => memory_space_6_lc_req(2 downto 2),
      memory_space_6_lc_ack => memory_space_6_lc_ack(2 downto 2),
      memory_space_6_lc_data => memory_space_6_lc_data(47 downto 32),
      memory_space_6_lc_tag => memory_space_6_lc_tag(2 downto 2),
      memory_space_7_lr_req => memory_space_7_lr_req(2 downto 2),
      memory_space_7_lr_ack => memory_space_7_lr_ack(2 downto 2),
      memory_space_7_lr_addr => memory_space_7_lr_addr(2 downto 2),
      memory_space_7_lr_tag => memory_space_7_lr_tag(59 downto 40),
      memory_space_7_lc_req => memory_space_7_lc_req(2 downto 2),
      memory_space_7_lc_ack => memory_space_7_lc_ack(2 downto 2),
      memory_space_7_lc_data => memory_space_7_lc_data(47 downto 32),
      memory_space_7_lc_tag => memory_space_7_lc_tag(5 downto 4),
      memory_space_5_sr_req => memory_space_5_sr_req(2 downto 2),
      memory_space_5_sr_ack => memory_space_5_sr_ack(2 downto 2),
      memory_space_5_sr_addr => memory_space_5_sr_addr(41 downto 28),
      memory_space_5_sr_data => memory_space_5_sr_data(191 downto 128),
      memory_space_5_sr_tag => memory_space_5_sr_tag(56 downto 38),
      memory_space_5_sc_req => memory_space_5_sc_req(2 downto 2),
      memory_space_5_sc_ack => memory_space_5_sc_ack(2 downto 2),
      memory_space_5_sc_tag => memory_space_5_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 7),
      memory_space_0_lr_tag => memory_space_0_lr_tag(41 downto 21),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 32),
      memory_space_0_lc_tag => memory_space_0_lc_tag(5 downto 3),
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 7),
      memory_space_1_lr_tag => memory_space_1_lr_tag(41 downto 21),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 32),
      memory_space_1_lc_tag => memory_space_1_lc_tag(5 downto 3),
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 1),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 1),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 7),
      memory_space_2_lr_tag => memory_space_2_lr_tag(39 downto 20),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 1),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 1),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 32),
      memory_space_2_lc_tag => memory_space_2_lc_tag(3 downto 2),
      memory_space_3_lr_req => memory_space_3_lr_req(1 downto 1),
      memory_space_3_lr_ack => memory_space_3_lr_ack(1 downto 1),
      memory_space_3_lr_addr => memory_space_3_lr_addr(27 downto 14),
      memory_space_3_lr_tag => memory_space_3_lr_tag(37 downto 19),
      memory_space_3_lc_req => memory_space_3_lc_req(1 downto 1),
      memory_space_3_lc_ack => memory_space_3_lc_ack(1 downto 1),
      memory_space_3_lc_data => memory_space_3_lc_data(127 downto 64),
      memory_space_3_lc_tag => memory_space_3_lc_tag(1 downto 1),
      memory_space_6_lr_req => memory_space_6_lr_req(1 downto 1),
      memory_space_6_lr_ack => memory_space_6_lr_ack(1 downto 1),
      memory_space_6_lr_addr => memory_space_6_lr_addr(1 downto 1),
      memory_space_6_lr_tag => memory_space_6_lr_tag(37 downto 19),
      memory_space_6_lc_req => memory_space_6_lc_req(1 downto 1),
      memory_space_6_lc_ack => memory_space_6_lc_ack(1 downto 1),
      memory_space_6_lc_data => memory_space_6_lc_data(31 downto 16),
      memory_space_6_lc_tag => memory_space_6_lc_tag(1 downto 1),
      memory_space_7_lr_req => memory_space_7_lr_req(1 downto 1),
      memory_space_7_lr_ack => memory_space_7_lr_ack(1 downto 1),
      memory_space_7_lr_addr => memory_space_7_lr_addr(1 downto 1),
      memory_space_7_lr_tag => memory_space_7_lr_tag(39 downto 20),
      memory_space_7_lc_req => memory_space_7_lc_req(1 downto 1),
      memory_space_7_lc_ack => memory_space_7_lc_ack(1 downto 1),
      memory_space_7_lc_data => memory_space_7_lc_data(31 downto 16),
      memory_space_7_lc_tag => memory_space_7_lc_tag(3 downto 2),
      memory_space_5_sr_req => memory_space_5_sr_req(1 downto 1),
      memory_space_5_sr_ack => memory_space_5_sr_ack(1 downto 1),
      memory_space_5_sr_addr => memory_space_5_sr_addr(27 downto 14),
      memory_space_5_sr_data => memory_space_5_sr_data(127 downto 64),
      memory_space_5_sr_tag => memory_space_5_sr_tag(37 downto 19),
      memory_space_5_sc_req => memory_space_5_sc_req(1 downto 1),
      memory_space_5_sc_ack => memory_space_5_sc_ack(1 downto 1),
      memory_space_5_sc_tag => memory_space_5_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(6 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(20 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(6 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(20 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(6 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(19 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(0 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(18 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(15 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(0 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(19 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(15 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(1 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(13 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(63 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(18 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(4 downto 4),
      memory_space_2_lr_ack => memory_space_2_lr_ack(4 downto 4),
      memory_space_2_lr_addr => memory_space_2_lr_addr(34 downto 28),
      memory_space_2_lr_tag => memory_space_2_lr_tag(99 downto 80),
      memory_space_2_lc_req => memory_space_2_lc_req(4 downto 4),
      memory_space_2_lc_ack => memory_space_2_lc_ack(4 downto 4),
      memory_space_2_lc_data => memory_space_2_lc_data(159 downto 128),
      memory_space_2_lc_tag => memory_space_2_lc_tag(9 downto 8),
      memory_space_5_lr_req => memory_space_5_lr_req(0 downto 0),
      memory_space_5_lr_ack => memory_space_5_lr_ack(0 downto 0),
      memory_space_5_lr_addr => memory_space_5_lr_addr(13 downto 0),
      memory_space_5_lr_tag => memory_space_5_lr_tag(18 downto 0),
      memory_space_5_lc_req => memory_space_5_lc_req(0 downto 0),
      memory_space_5_lc_ack => memory_space_5_lc_ack(0 downto 0),
      memory_space_5_lc_data => memory_space_5_lc_data(63 downto 0),
      memory_space_5_lc_tag => memory_space_5_lc_tag(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module testConfigure
  testConfigure_out_args <= testConfigure_ret_val_x_x ;
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      return_data =>testConfigure_return_data,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      return_mdata => testConfigure_out_args,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => testConfigure_ret_val_x_x,
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(4 downto 4),
      memory_space_0_lr_ack => memory_space_0_lr_ack(4 downto 4),
      memory_space_0_lr_addr => memory_space_0_lr_addr(34 downto 28),
      memory_space_0_lr_tag => memory_space_0_lr_tag(104 downto 84),
      memory_space_0_lc_req => memory_space_0_lc_req(4 downto 4),
      memory_space_0_lc_ack => memory_space_0_lc_ack(4 downto 4),
      memory_space_0_lc_data => memory_space_0_lc_data(159 downto 128),
      memory_space_0_lc_tag => memory_space_0_lc_tag(14 downto 12),
      memory_space_1_lr_req => memory_space_1_lr_req(4 downto 4),
      memory_space_1_lr_ack => memory_space_1_lr_ack(4 downto 4),
      memory_space_1_lr_addr => memory_space_1_lr_addr(34 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(104 downto 84),
      memory_space_1_lc_req => memory_space_1_lc_req(4 downto 4),
      memory_space_1_lc_ack => memory_space_1_lc_ack(4 downto 4),
      memory_space_1_lc_data => memory_space_1_lc_data(159 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(14 downto 12),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(6 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(20 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(6 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(20 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(2 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(6 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(19 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(10 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(63 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(0 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(0 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(15 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(18 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(0 downto 0),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(15 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(19 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(1 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_4: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_loads => 1,
      num_stores => 4,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
