-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity concat is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    Concat_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    Concat_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Concat_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Concat_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity concat;
architecture concat_arch of concat is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal concat_CP_34_start: Boolean;
  signal concat_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_755_call_req_1 : boolean;
  signal if_stmt_744_branch_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_610_inst_ack_1 : boolean;
  signal call_stmt_755_call_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_610_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_646_inst_ack_1 : boolean;
  signal type_cast_614_inst_ack_1 : boolean;
  signal type_cast_614_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_51_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_51_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_610_inst_ack_0 : boolean;
  signal array_obj_ref_593_index_offset_ack_1 : boolean;
  signal array_obj_ref_593_index_offset_req_1 : boolean;
  signal type_cast_614_inst_ack_0 : boolean;
  signal type_cast_614_inst_req_0 : boolean;
  signal array_obj_ref_593_index_offset_ack_0 : boolean;
  signal type_cast_956_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_25_inst_req_0 : boolean;
  signal type_cast_668_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_25_inst_ack_0 : boolean;
  signal type_cast_686_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_25_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_25_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_646_inst_req_1 : boolean;
  signal type_cast_30_inst_req_0 : boolean;
  signal type_cast_668_inst_req_1 : boolean;
  signal type_cast_30_inst_ack_0 : boolean;
  signal type_cast_30_inst_req_1 : boolean;
  signal type_cast_30_inst_ack_1 : boolean;
  signal call_stmt_755_call_req_0 : boolean;
  signal type_cast_686_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_39_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_39_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_39_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_39_inst_ack_1 : boolean;
  signal array_obj_ref_845_index_offset_req_0 : boolean;
  signal type_cast_43_inst_req_0 : boolean;
  signal type_cast_43_inst_ack_0 : boolean;
  signal type_cast_43_inst_req_1 : boolean;
  signal type_cast_43_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_51_inst_req_0 : boolean;
  signal type_cast_668_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_51_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_610_inst_req_0 : boolean;
  signal type_cast_986_inst_ack_0 : boolean;
  signal call_stmt_917_call_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1011_inst_ack_1 : boolean;
  signal type_cast_143_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_664_inst_req_1 : boolean;
  signal type_cast_143_inst_ack_0 : boolean;
  signal type_cast_143_inst_req_1 : boolean;
  signal type_cast_143_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_646_inst_ack_0 : boolean;
  signal type_cast_55_inst_req_0 : boolean;
  signal type_cast_668_inst_req_0 : boolean;
  signal type_cast_55_inst_ack_0 : boolean;
  signal type_cast_55_inst_req_1 : boolean;
  signal type_cast_956_inst_ack_1 : boolean;
  signal type_cast_55_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_64_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_64_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_64_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_64_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_646_inst_req_0 : boolean;
  signal type_cast_68_inst_req_0 : boolean;
  signal phi_stmt_581_ack_0 : boolean;
  signal type_cast_68_inst_ack_0 : boolean;
  signal type_cast_936_inst_req_1 : boolean;
  signal type_cast_68_inst_req_1 : boolean;
  signal type_cast_68_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_76_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_76_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_76_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_76_inst_ack_1 : boolean;
  signal SUB_u32_u32_903_inst_ack_1 : boolean;
  signal do_while_stmt_784_branch_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_718_inst_ack_1 : boolean;
  signal type_cast_80_inst_req_0 : boolean;
  signal type_cast_80_inst_ack_0 : boolean;
  signal type_cast_80_inst_req_1 : boolean;
  signal type_cast_80_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_89_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_89_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_89_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_89_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_718_inst_req_1 : boolean;
  signal type_cast_93_inst_req_0 : boolean;
  signal type_cast_93_inst_ack_0 : boolean;
  signal type_cast_93_inst_req_1 : boolean;
  signal type_cast_93_inst_ack_1 : boolean;
  signal do_while_stmt_784_branch_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_700_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_101_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_101_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_101_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_101_inst_ack_1 : boolean;
  signal SUB_u32_u32_903_inst_ack_0 : boolean;
  signal if_stmt_744_branch_ack_0 : boolean;
  signal do_while_stmt_784_branch_ack_1 : boolean;
  signal array_obj_ref_845_index_offset_ack_0 : boolean;
  signal type_cast_105_inst_req_0 : boolean;
  signal type_cast_105_inst_ack_0 : boolean;
  signal type_cast_105_inst_req_1 : boolean;
  signal type_cast_105_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_700_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_114_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_114_inst_ack_0 : boolean;
  signal type_cast_601_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1008_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_114_inst_req_1 : boolean;
  signal call_stmt_917_call_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_114_inst_ack_1 : boolean;
  signal W_cmp_844_delayed_12_0_851_inst_req_0 : boolean;
  signal type_cast_118_inst_req_0 : boolean;
  signal type_cast_118_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_718_inst_ack_0 : boolean;
  signal type_cast_118_inst_req_1 : boolean;
  signal type_cast_118_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_700_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_126_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_126_inst_ack_0 : boolean;
  signal type_cast_601_inst_req_1 : boolean;
  signal SUB_u32_u32_903_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_126_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_126_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1011_inst_req_1 : boolean;
  signal type_cast_936_inst_ack_1 : boolean;
  signal type_cast_130_inst_req_0 : boolean;
  signal type_cast_130_inst_ack_0 : boolean;
  signal array_obj_ref_593_index_offset_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_718_inst_req_0 : boolean;
  signal type_cast_130_inst_req_1 : boolean;
  signal type_cast_130_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_700_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_139_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_664_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_139_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_139_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_139_inst_ack_1 : boolean;
  signal array_obj_ref_386_index_offset_ack_0 : boolean;
  signal array_obj_ref_386_index_offset_req_1 : boolean;
  signal array_obj_ref_386_index_offset_ack_1 : boolean;
  signal MUX_859_inst_ack_0 : boolean;
  signal type_cast_922_inst_req_0 : boolean;
  signal addr_of_387_final_reg_req_0 : boolean;
  signal addr_of_387_final_reg_ack_0 : boolean;
  signal addr_of_387_final_reg_req_1 : boolean;
  signal addr_of_387_final_reg_ack_1 : boolean;
  signal type_cast_946_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_151_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_151_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_151_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_151_inst_ack_1 : boolean;
  signal type_cast_956_inst_req_0 : boolean;
  signal type_cast_722_inst_ack_1 : boolean;
  signal type_cast_722_inst_req_1 : boolean;
  signal type_cast_155_inst_req_0 : boolean;
  signal type_cast_155_inst_ack_0 : boolean;
  signal type_cast_155_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_664_inst_ack_0 : boolean;
  signal type_cast_155_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_682_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_164_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_164_inst_ack_0 : boolean;
  signal type_cast_601_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_164_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_664_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_164_inst_ack_1 : boolean;
  signal ptr_deref_730_store_0_ack_1 : boolean;
  signal if_stmt_744_branch_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_682_inst_req_1 : boolean;
  signal type_cast_168_inst_req_0 : boolean;
  signal type_cast_168_inst_ack_0 : boolean;
  signal type_cast_168_inst_req_1 : boolean;
  signal type_cast_168_inst_ack_1 : boolean;
  signal W_cmp_844_delayed_12_0_851_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_176_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_176_inst_ack_0 : boolean;
  signal type_cast_601_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_176_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_176_inst_ack_1 : boolean;
  signal ptr_deref_730_store_0_req_1 : boolean;
  signal type_cast_722_inst_ack_0 : boolean;
  signal call_stmt_917_call_ack_1 : boolean;
  signal type_cast_722_inst_req_0 : boolean;
  signal type_cast_181_inst_req_0 : boolean;
  signal type_cast_181_inst_ack_0 : boolean;
  signal type_cast_181_inst_req_1 : boolean;
  signal type_cast_181_inst_ack_1 : boolean;
  signal W_cmp_844_delayed_12_0_851_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_682_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_190_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_190_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_190_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_190_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1020_inst_ack_1 : boolean;
  signal type_cast_194_inst_req_0 : boolean;
  signal type_cast_194_inst_ack_0 : boolean;
  signal type_cast_194_inst_req_1 : boolean;
  signal type_cast_194_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_682_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_202_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_202_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_202_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_202_inst_ack_1 : boolean;
  signal call_stmt_755_call_ack_1 : boolean;
  signal type_cast_632_inst_ack_1 : boolean;
  signal type_cast_632_inst_req_1 : boolean;
  signal addr_of_846_final_reg_req_0 : boolean;
  signal type_cast_206_inst_req_0 : boolean;
  signal type_cast_206_inst_ack_0 : boolean;
  signal type_cast_206_inst_req_1 : boolean;
  signal type_cast_206_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_215_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_215_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_597_inst_ack_1 : boolean;
  signal type_cast_936_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_215_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_215_inst_ack_1 : boolean;
  signal type_cast_632_inst_ack_0 : boolean;
  signal type_cast_219_inst_req_0 : boolean;
  signal type_cast_219_inst_ack_0 : boolean;
  signal type_cast_219_inst_req_1 : boolean;
  signal type_cast_219_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_597_inst_req_1 : boolean;
  signal type_cast_936_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_227_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_227_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_227_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_227_inst_ack_1 : boolean;
  signal type_cast_632_inst_req_0 : boolean;
  signal type_cast_650_inst_ack_1 : boolean;
  signal type_cast_231_inst_req_0 : boolean;
  signal call_stmt_917_call_ack_0 : boolean;
  signal type_cast_231_inst_ack_0 : boolean;
  signal type_cast_231_inst_req_1 : boolean;
  signal type_cast_650_inst_req_1 : boolean;
  signal type_cast_231_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_597_inst_ack_0 : boolean;
  signal type_cast_686_inst_ack_1 : boolean;
  signal type_cast_956_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_240_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_240_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_597_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_240_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_240_inst_ack_1 : boolean;
  signal type_cast_244_inst_req_0 : boolean;
  signal type_cast_244_inst_ack_0 : boolean;
  signal type_cast_244_inst_req_1 : boolean;
  signal type_cast_650_inst_ack_0 : boolean;
  signal type_cast_244_inst_ack_1 : boolean;
  signal W_cmp_844_delayed_12_0_851_inst_ack_0 : boolean;
  signal type_cast_258_inst_req_0 : boolean;
  signal type_cast_650_inst_req_0 : boolean;
  signal type_cast_258_inst_ack_0 : boolean;
  signal type_cast_704_inst_ack_1 : boolean;
  signal type_cast_258_inst_req_1 : boolean;
  signal type_cast_258_inst_ack_1 : boolean;
  signal type_cast_262_inst_req_0 : boolean;
  signal type_cast_262_inst_ack_0 : boolean;
  signal type_cast_704_inst_req_1 : boolean;
  signal type_cast_262_inst_req_1 : boolean;
  signal type_cast_262_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_628_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_628_inst_req_1 : boolean;
  signal type_cast_276_inst_req_0 : boolean;
  signal type_cast_276_inst_ack_0 : boolean;
  signal type_cast_276_inst_req_1 : boolean;
  signal type_cast_276_inst_ack_1 : boolean;
  signal addr_of_594_final_reg_ack_1 : boolean;
  signal addr_of_594_final_reg_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_628_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_628_inst_req_0 : boolean;
  signal type_cast_280_inst_req_0 : boolean;
  signal type_cast_280_inst_ack_0 : boolean;
  signal type_cast_280_inst_req_1 : boolean;
  signal type_cast_280_inst_ack_1 : boolean;
  signal ptr_deref_730_store_0_ack_0 : boolean;
  signal ptr_deref_730_store_0_req_0 : boolean;
  signal type_cast_686_inst_req_1 : boolean;
  signal type_cast_704_inst_ack_0 : boolean;
  signal addr_of_594_final_reg_ack_0 : boolean;
  signal if_stmt_315_branch_req_0 : boolean;
  signal if_stmt_315_branch_ack_1 : boolean;
  signal if_stmt_315_branch_ack_0 : boolean;
  signal type_cast_704_inst_req_0 : boolean;
  signal addr_of_594_final_reg_req_0 : boolean;
  signal if_stmt_330_branch_req_0 : boolean;
  signal addr_of_846_final_reg_ack_0 : boolean;
  signal if_stmt_330_branch_ack_1 : boolean;
  signal if_stmt_330_branch_ack_0 : boolean;
  signal type_cast_357_inst_req_0 : boolean;
  signal type_cast_357_inst_ack_0 : boolean;
  signal type_cast_357_inst_req_1 : boolean;
  signal type_cast_357_inst_ack_1 : boolean;
  signal type_cast_946_inst_req_0 : boolean;
  signal MUX_859_inst_req_0 : boolean;
  signal array_obj_ref_386_index_offset_req_0 : boolean;
  signal type_cast_922_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_390_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_390_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_390_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_390_inst_ack_1 : boolean;
  signal phi_stmt_374_req_1 : boolean;
  signal addr_of_846_final_reg_req_1 : boolean;
  signal type_cast_394_inst_req_0 : boolean;
  signal type_cast_394_inst_ack_0 : boolean;
  signal type_cast_394_inst_req_1 : boolean;
  signal type_cast_394_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_403_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_403_inst_ack_0 : boolean;
  signal MUX_859_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_403_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_403_inst_ack_1 : boolean;
  signal type_cast_922_inst_req_1 : boolean;
  signal type_cast_922_inst_ack_1 : boolean;
  signal type_cast_407_inst_req_0 : boolean;
  signal type_cast_407_inst_ack_0 : boolean;
  signal type_cast_407_inst_req_1 : boolean;
  signal type_cast_407_inst_ack_1 : boolean;
  signal type_cast_380_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_421_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_421_inst_ack_0 : boolean;
  signal MUX_859_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_421_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_421_inst_ack_1 : boolean;
  signal array_obj_ref_845_index_offset_req_1 : boolean;
  signal type_cast_425_inst_req_0 : boolean;
  signal type_cast_425_inst_ack_0 : boolean;
  signal type_cast_425_inst_req_1 : boolean;
  signal type_cast_425_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_439_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_439_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_439_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_439_inst_ack_1 : boolean;
  signal addr_of_846_final_reg_ack_1 : boolean;
  signal type_cast_927_inst_req_0 : boolean;
  signal type_cast_443_inst_req_0 : boolean;
  signal type_cast_443_inst_ack_0 : boolean;
  signal type_cast_443_inst_req_1 : boolean;
  signal array_obj_ref_845_index_offset_ack_1 : boolean;
  signal type_cast_443_inst_ack_1 : boolean;
  signal type_cast_986_inst_req_0 : boolean;
  signal type_cast_927_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_457_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_457_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_457_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_457_inst_ack_1 : boolean;
  signal type_cast_461_inst_req_0 : boolean;
  signal type_cast_461_inst_ack_0 : boolean;
  signal type_cast_461_inst_req_1 : boolean;
  signal type_cast_461_inst_ack_1 : boolean;
  signal type_cast_927_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_475_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_475_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_475_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_475_inst_ack_1 : boolean;
  signal type_cast_479_inst_req_0 : boolean;
  signal type_cast_479_inst_ack_0 : boolean;
  signal type_cast_479_inst_req_1 : boolean;
  signal type_cast_479_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_493_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_493_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_493_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_493_inst_ack_1 : boolean;
  signal type_cast_497_inst_req_0 : boolean;
  signal type_cast_497_inst_ack_0 : boolean;
  signal type_cast_497_inst_req_1 : boolean;
  signal type_cast_497_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_511_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_511_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_511_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_511_inst_ack_1 : boolean;
  signal type_cast_515_inst_req_0 : boolean;
  signal type_cast_515_inst_ack_0 : boolean;
  signal type_cast_515_inst_req_1 : boolean;
  signal type_cast_515_inst_ack_1 : boolean;
  signal ptr_deref_523_store_0_req_0 : boolean;
  signal ptr_deref_523_store_0_ack_0 : boolean;
  signal ptr_deref_523_store_0_req_1 : boolean;
  signal ptr_deref_523_store_0_ack_1 : boolean;
  signal if_stmt_537_branch_req_0 : boolean;
  signal if_stmt_537_branch_ack_1 : boolean;
  signal if_stmt_537_branch_ack_0 : boolean;
  signal type_cast_564_inst_req_0 : boolean;
  signal type_cast_564_inst_ack_0 : boolean;
  signal type_cast_564_inst_req_1 : boolean;
  signal type_cast_564_inst_ack_1 : boolean;
  signal type_cast_996_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1014_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1014_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1008_inst_req_1 : boolean;
  signal phi_stmt_786_req_1 : boolean;
  signal phi_stmt_786_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1008_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1023_inst_req_1 : boolean;
  signal phi_stmt_786_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1008_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1011_inst_ack_0 : boolean;
  signal type_cast_976_inst_ack_1 : boolean;
  signal type_cast_976_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1011_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1014_inst_ack_0 : boolean;
  signal type_cast_976_inst_ack_0 : boolean;
  signal type_cast_976_inst_req_0 : boolean;
  signal next_add_out_899_789_buf_req_0 : boolean;
  signal next_add_out_899_789_buf_ack_0 : boolean;
  signal SUB_u32_u32_903_inst_req_0 : boolean;
  signal type_cast_587_inst_ack_1 : boolean;
  signal next_add_out_899_789_buf_req_1 : boolean;
  signal next_add_out_899_789_buf_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1014_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1020_inst_req_1 : boolean;
  signal type_cast_996_inst_req_1 : boolean;
  signal phi_stmt_790_req_1 : boolean;
  signal phi_stmt_790_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1017_inst_ack_1 : boolean;
  signal phi_stmt_790_ack_0 : boolean;
  signal phi_stmt_581_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1020_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1017_inst_req_1 : boolean;
  signal SUB_u16_u16_864_inst_ack_1 : boolean;
  signal next_add_inp1_886_793_buf_req_0 : boolean;
  signal next_add_inp1_886_793_buf_ack_0 : boolean;
  signal SUB_u16_u16_864_inst_req_1 : boolean;
  signal next_add_inp1_886_793_buf_req_1 : boolean;
  signal next_add_inp1_886_793_buf_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1020_inst_req_0 : boolean;
  signal SUB_u16_u16_864_inst_ack_0 : boolean;
  signal SUB_u16_u16_864_inst_req_0 : boolean;
  signal phi_stmt_581_req_1 : boolean;
  signal type_cast_380_inst_req_1 : boolean;
  signal phi_stmt_794_req_1 : boolean;
  signal type_cast_1006_inst_ack_1 : boolean;
  signal phi_stmt_794_req_0 : boolean;
  signal type_cast_1006_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1023_inst_ack_0 : boolean;
  signal type_cast_996_inst_ack_0 : boolean;
  signal phi_stmt_794_ack_0 : boolean;
  signal type_cast_986_inst_ack_1 : boolean;
  signal type_cast_1006_inst_ack_0 : boolean;
  signal type_cast_986_inst_req_1 : boolean;
  signal type_cast_1083_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1017_inst_ack_0 : boolean;
  signal next_add_inp2_894_797_buf_req_0 : boolean;
  signal next_add_inp2_894_797_buf_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1017_inst_req_0 : boolean;
  signal next_add_inp2_894_797_buf_req_1 : boolean;
  signal next_add_inp2_894_797_buf_ack_1 : boolean;
  signal ptr_deref_855_store_0_ack_1 : boolean;
  signal type_cast_1006_inst_req_0 : boolean;
  signal phi_stmt_798_req_1 : boolean;
  signal phi_stmt_1077_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1023_inst_req_0 : boolean;
  signal phi_stmt_798_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1023_inst_ack_1 : boolean;
  signal type_cast_996_inst_req_0 : boolean;
  signal phi_stmt_798_ack_0 : boolean;
  signal type_cast_966_inst_ack_1 : boolean;
  signal type_cast_927_inst_ack_1 : boolean;
  signal ptr_deref_855_store_0_req_1 : boolean;
  signal type_cast_966_inst_req_1 : boolean;
  signal next_count_inp1_878_801_buf_req_0 : boolean;
  signal next_count_inp1_878_801_buf_ack_0 : boolean;
  signal next_count_inp1_878_801_buf_req_1 : boolean;
  signal next_count_inp1_878_801_buf_ack_1 : boolean;
  signal ptr_deref_855_store_0_ack_0 : boolean;
  signal ptr_deref_855_store_0_req_0 : boolean;
  signal W_ov_842_delayed_7_0_848_inst_ack_1 : boolean;
  signal array_obj_ref_813_index_offset_req_0 : boolean;
  signal array_obj_ref_813_index_offset_ack_0 : boolean;
  signal W_ov_842_delayed_7_0_848_inst_req_1 : boolean;
  signal array_obj_ref_813_index_offset_req_1 : boolean;
  signal array_obj_ref_813_index_offset_ack_1 : boolean;
  signal addr_of_814_final_reg_req_0 : boolean;
  signal addr_of_814_final_reg_ack_0 : boolean;
  signal addr_of_814_final_reg_req_1 : boolean;
  signal type_cast_946_inst_ack_1 : boolean;
  signal addr_of_814_final_reg_ack_1 : boolean;
  signal W_ov_842_delayed_7_0_848_inst_ack_0 : boolean;
  signal type_cast_966_inst_ack_0 : boolean;
  signal W_ov_842_delayed_7_0_848_inst_req_0 : boolean;
  signal W_cmp_816_delayed_6_0_816_inst_req_0 : boolean;
  signal type_cast_946_inst_req_1 : boolean;
  signal W_cmp_816_delayed_6_0_816_inst_ack_0 : boolean;
  signal W_cmp_816_delayed_6_0_816_inst_req_1 : boolean;
  signal W_cmp_816_delayed_6_0_816_inst_ack_1 : boolean;
  signal type_cast_966_inst_req_0 : boolean;
  signal phi_stmt_374_req_0 : boolean;
  signal type_cast_1083_inst_ack_0 : boolean;
  signal ptr_deref_822_load_0_req_0 : boolean;
  signal ptr_deref_822_load_0_ack_0 : boolean;
  signal ptr_deref_822_load_0_req_1 : boolean;
  signal ptr_deref_822_load_0_ack_1 : boolean;
  signal type_cast_1083_inst_req_1 : boolean;
  signal array_obj_ref_829_index_offset_req_0 : boolean;
  signal array_obj_ref_829_index_offset_ack_0 : boolean;
  signal type_cast_1083_inst_ack_1 : boolean;
  signal array_obj_ref_829_index_offset_req_1 : boolean;
  signal array_obj_ref_829_index_offset_ack_1 : boolean;
  signal phi_stmt_1077_req_1 : boolean;
  signal addr_of_830_final_reg_req_0 : boolean;
  signal addr_of_830_final_reg_ack_0 : boolean;
  signal addr_of_830_final_reg_req_1 : boolean;
  signal addr_of_830_final_reg_ack_1 : boolean;
  signal W_cmp_829_delayed_6_0_832_inst_req_0 : boolean;
  signal W_cmp_829_delayed_6_0_832_inst_ack_0 : boolean;
  signal W_cmp_829_delayed_6_0_832_inst_req_1 : boolean;
  signal W_cmp_829_delayed_6_0_832_inst_ack_1 : boolean;
  signal ptr_deref_838_load_0_req_0 : boolean;
  signal ptr_deref_838_load_0_ack_0 : boolean;
  signal ptr_deref_838_load_0_req_1 : boolean;
  signal ptr_deref_838_load_0_ack_1 : boolean;
  signal type_cast_380_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1026_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1026_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1026_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1026_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1029_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1029_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1029_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1029_inst_ack_1 : boolean;
  signal type_cast_587_inst_req_1 : boolean;
  signal type_cast_380_inst_req_0 : boolean;
  signal if_stmt_1039_branch_req_0 : boolean;
  signal if_stmt_1039_branch_ack_1 : boolean;
  signal if_stmt_1039_branch_ack_0 : boolean;
  signal type_cast_1060_inst_req_0 : boolean;
  signal type_cast_1060_inst_ack_0 : boolean;
  signal type_cast_1060_inst_req_1 : boolean;
  signal type_cast_1060_inst_ack_1 : boolean;
  signal array_obj_ref_1089_index_offset_req_0 : boolean;
  signal array_obj_ref_1089_index_offset_ack_0 : boolean;
  signal array_obj_ref_1089_index_offset_req_1 : boolean;
  signal array_obj_ref_1089_index_offset_ack_1 : boolean;
  signal addr_of_1090_final_reg_req_0 : boolean;
  signal addr_of_1090_final_reg_ack_0 : boolean;
  signal addr_of_1090_final_reg_req_1 : boolean;
  signal addr_of_1090_final_reg_ack_1 : boolean;
  signal type_cast_587_inst_ack_0 : boolean;
  signal type_cast_587_inst_req_0 : boolean;
  signal ptr_deref_1094_load_0_req_0 : boolean;
  signal ptr_deref_1094_load_0_ack_0 : boolean;
  signal ptr_deref_1094_load_0_req_1 : boolean;
  signal ptr_deref_1094_load_0_ack_1 : boolean;
  signal type_cast_1098_inst_req_0 : boolean;
  signal type_cast_1098_inst_ack_0 : boolean;
  signal type_cast_1098_inst_req_1 : boolean;
  signal type_cast_1098_inst_ack_1 : boolean;
  signal type_cast_1108_inst_req_0 : boolean;
  signal type_cast_1108_inst_ack_0 : boolean;
  signal type_cast_1108_inst_req_1 : boolean;
  signal type_cast_1108_inst_ack_1 : boolean;
  signal type_cast_1118_inst_req_0 : boolean;
  signal type_cast_1118_inst_ack_0 : boolean;
  signal type_cast_1118_inst_req_1 : boolean;
  signal type_cast_1118_inst_ack_1 : boolean;
  signal type_cast_1128_inst_req_0 : boolean;
  signal type_cast_1128_inst_ack_0 : boolean;
  signal type_cast_1128_inst_req_1 : boolean;
  signal type_cast_1128_inst_ack_1 : boolean;
  signal type_cast_1138_inst_req_0 : boolean;
  signal type_cast_1138_inst_ack_0 : boolean;
  signal type_cast_1138_inst_req_1 : boolean;
  signal type_cast_1138_inst_ack_1 : boolean;
  signal type_cast_1148_inst_req_0 : boolean;
  signal type_cast_1148_inst_ack_0 : boolean;
  signal type_cast_1148_inst_req_1 : boolean;
  signal type_cast_1148_inst_ack_1 : boolean;
  signal type_cast_1158_inst_req_0 : boolean;
  signal type_cast_1158_inst_ack_0 : boolean;
  signal type_cast_1158_inst_req_1 : boolean;
  signal type_cast_1158_inst_ack_1 : boolean;
  signal type_cast_1168_inst_req_0 : boolean;
  signal type_cast_1168_inst_ack_0 : boolean;
  signal type_cast_1168_inst_req_1 : boolean;
  signal type_cast_1168_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1170_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1170_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1170_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1170_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1173_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1173_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1173_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1173_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1176_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1176_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1176_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1176_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1179_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1179_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1179_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1179_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1182_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1182_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1182_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1182_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1185_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1185_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1185_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1185_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1188_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1188_inst_ack_0 : boolean;
  signal phi_stmt_374_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1188_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1188_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1191_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1191_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1191_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1191_inst_ack_1 : boolean;
  signal if_stmt_1205_branch_req_0 : boolean;
  signal if_stmt_1205_branch_ack_1 : boolean;
  signal phi_stmt_1077_ack_0 : boolean;
  signal if_stmt_1205_branch_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "concat_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  concat_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "concat_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= concat_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= concat_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= concat_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  concat_CP_34: Block -- control-path 
    signal concat_CP_34_elements: BooleanArray(459 downto 0);
    -- 
  begin -- 
    concat_CP_34_elements(0) <= concat_CP_34_start;
    concat_CP_34_symbol <= concat_CP_34_elements(459);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	82 
    -- CP-element group 0: 	53 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	61 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	73 
    -- CP-element group 0: 	76 
    -- CP-element group 0: 	79 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	17 
    -- CP-element group 0:  members (74) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_23/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/branch_block_stmt_23__entry__
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314__entry__
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_25_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_25_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_25_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_30_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_30_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_30_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_43_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_43_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_43_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_143_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_143_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_143_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_55_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_55_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_55_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_68_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_68_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_68_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_80_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_80_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_80_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_93_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_93_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_93_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_105_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_105_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_105_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_118_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_118_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_118_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_130_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_130_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_130_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_155_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_155_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_155_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_168_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_168_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_168_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_181_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_181_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_181_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_194_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_194_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_194_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_206_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_206_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_206_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_219_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_219_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_219_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_231_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_231_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_231_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_244_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_244_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_244_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_258_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_258_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_258_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_262_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_262_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_262_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_276_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_276_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_276_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_280_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_280_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_280_Update/cr
      -- 
    rr_116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => RPIPE_Concat_input_pipe_25_inst_req_0); -- 
    cr_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_30_inst_req_1); -- 
    cr_163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_43_inst_req_1); -- 
    cr_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_143_inst_req_1); -- 
    cr_191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_55_inst_req_1); -- 
    cr_219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_68_inst_req_1); -- 
    cr_247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_80_inst_req_1); -- 
    cr_275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_93_inst_req_1); -- 
    cr_303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_105_inst_req_1); -- 
    cr_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_118_inst_req_1); -- 
    cr_359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_130_inst_req_1); -- 
    cr_415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_155_inst_req_1); -- 
    cr_443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_168_inst_req_1); -- 
    cr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_181_inst_req_1); -- 
    cr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_194_inst_req_1); -- 
    cr_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_206_inst_req_1); -- 
    cr_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_219_inst_req_1); -- 
    cr_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_231_inst_req_1); -- 
    cr_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_244_inst_req_1); -- 
    cr_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_258_inst_req_1); -- 
    cr_639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_262_inst_req_1); -- 
    cr_653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_276_inst_req_1); -- 
    cr_667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_280_inst_req_1); -- 
    -- CP-element group 1:  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	333 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	334 
    -- CP-element group 1: 	335 
    -- CP-element group 1: 	336 
    -- CP-element group 1: 	337 
    -- CP-element group 1: 	339 
    -- CP-element group 1: 	342 
    -- CP-element group 1: 	345 
    -- CP-element group 1: 	348 
    -- CP-element group 1: 	351 
    -- CP-element group 1: 	354 
    -- CP-element group 1: 	357 
    -- CP-element group 1: 	360 
    -- CP-element group 1: 	363 
    -- CP-element group 1:  members (42) 
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/call_stmt_917_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/do_while_stmt_784__exit__
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031__entry__
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_956_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/call_stmt_917_Update/ccr
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_956_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_936_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/call_stmt_917_Sample/crr
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/call_stmt_917_update_start_
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_922_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_946_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/call_stmt_917_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_936_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_922_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_922_update_start_
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_996_update_start_
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_986_update_start_
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/call_stmt_917_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_946_update_start_
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_922_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_966_update_start_
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_922_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_922_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_927_update_start_
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_927_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_927_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_976_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_976_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_936_update_start_
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_996_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_976_update_start_
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_996_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_1006_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_1006_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_986_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_1006_update_start_
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_966_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_986_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_966_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_956_update_start_
      -- CP-element group 1: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_946_Update/cr
      -- 
    cr_2125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => type_cast_956_inst_req_1); -- 
    ccr_2055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => call_stmt_917_call_req_1); -- 
    cr_2097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => type_cast_936_inst_req_1); -- 
    crr_2050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => call_stmt_917_call_req_0); -- 
    rr_2064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => type_cast_922_inst_req_0); -- 
    cr_2069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => type_cast_922_inst_req_1); -- 
    cr_2083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => type_cast_927_inst_req_1); -- 
    cr_2153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => type_cast_976_inst_req_1); -- 
    cr_2181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => type_cast_996_inst_req_1); -- 
    cr_2195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => type_cast_1006_inst_req_1); -- 
    cr_2167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => type_cast_986_inst_req_1); -- 
    cr_2139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => type_cast_966_inst_req_1); -- 
    cr_2111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => type_cast_946_inst_req_1); -- 
    concat_CP_34_elements(1) <= concat_CP_34_elements(333);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_25_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_25_update_start_
      -- CP-element group 2: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_25_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_25_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_25_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_25_Update/cr
      -- 
    ra_117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_25_inst_ack_0, ack => concat_CP_34_elements(2)); -- 
    cr_121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(2), ack => RPIPE_Concat_input_pipe_25_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_25_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_25_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_25_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_30_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_30_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_30_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_39_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_39_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_39_Sample/rr
      -- 
    ca_122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_25_inst_ack_1, ack => concat_CP_34_elements(3)); -- 
    rr_130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(3), ack => type_cast_30_inst_req_0); -- 
    rr_144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(3), ack => RPIPE_Concat_input_pipe_39_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_30_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_30_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_30_Sample/ra
      -- 
    ra_131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_30_inst_ack_0, ack => concat_CP_34_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	77 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_30_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_30_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_30_Update/ca
      -- 
    ca_136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_30_inst_ack_1, ack => concat_CP_34_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_39_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_39_update_start_
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_39_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_39_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_39_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_39_Update/cr
      -- 
    ra_145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_39_inst_ack_0, ack => concat_CP_34_elements(6)); -- 
    cr_149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(6), ack => RPIPE_Concat_input_pipe_39_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_39_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_39_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_39_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_43_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_43_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_43_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_51_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_51_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_51_Sample/rr
      -- 
    ca_150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_39_inst_ack_1, ack => concat_CP_34_elements(7)); -- 
    rr_158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(7), ack => type_cast_43_inst_req_0); -- 
    rr_172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(7), ack => RPIPE_Concat_input_pipe_51_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_43_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_43_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_43_Sample/ra
      -- 
    ra_159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_43_inst_ack_0, ack => concat_CP_34_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	77 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_43_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_43_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_43_Update/ca
      -- 
    ca_164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_43_inst_ack_1, ack => concat_CP_34_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_51_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_51_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_51_update_start_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_51_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_51_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_51_Update/$entry
      -- 
    ra_173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_51_inst_ack_0, ack => concat_CP_34_elements(10)); -- 
    cr_177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(10), ack => RPIPE_Concat_input_pipe_51_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_51_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_55_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_51_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_51_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_55_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_55_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_64_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_64_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_64_Sample/rr
      -- 
    ca_178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_51_inst_ack_1, ack => concat_CP_34_elements(11)); -- 
    rr_186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(11), ack => type_cast_55_inst_req_0); -- 
    rr_200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(11), ack => RPIPE_Concat_input_pipe_64_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_55_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_55_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_55_Sample/ra
      -- 
    ra_187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_55_inst_ack_0, ack => concat_CP_34_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	74 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_55_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_55_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_55_Update/ca
      -- 
    ca_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_55_inst_ack_1, ack => concat_CP_34_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_64_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_64_update_start_
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_64_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_64_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_64_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_64_Update/cr
      -- 
    ra_201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_64_inst_ack_0, ack => concat_CP_34_elements(14)); -- 
    cr_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(14), ack => RPIPE_Concat_input_pipe_64_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_64_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_64_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_64_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_68_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_68_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_68_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_76_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_76_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_76_Sample/rr
      -- 
    ca_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_64_inst_ack_1, ack => concat_CP_34_elements(15)); -- 
    rr_214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(15), ack => type_cast_68_inst_req_0); -- 
    rr_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(15), ack => RPIPE_Concat_input_pipe_76_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_68_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_68_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_68_Sample/ra
      -- 
    ra_215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_68_inst_ack_0, ack => concat_CP_34_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	74 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_68_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_68_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_68_Update/ca
      -- 
    ca_220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_68_inst_ack_1, ack => concat_CP_34_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_76_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_76_update_start_
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_76_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_76_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_76_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_76_Update/cr
      -- 
    ra_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_76_inst_ack_0, ack => concat_CP_34_elements(18)); -- 
    cr_233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(18), ack => RPIPE_Concat_input_pipe_76_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_76_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_76_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_76_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_80_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_80_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_80_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_89_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_89_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_89_Sample/rr
      -- 
    ca_234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_76_inst_ack_1, ack => concat_CP_34_elements(19)); -- 
    rr_242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(19), ack => type_cast_80_inst_req_0); -- 
    rr_256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(19), ack => RPIPE_Concat_input_pipe_89_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_80_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_80_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_80_Sample/ra
      -- 
    ra_243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_80_inst_ack_0, ack => concat_CP_34_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	74 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_80_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_80_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_80_Update/ca
      -- 
    ca_248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_80_inst_ack_1, ack => concat_CP_34_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_89_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_89_update_start_
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_89_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_89_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_89_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_89_Update/cr
      -- 
    ra_257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_89_inst_ack_0, ack => concat_CP_34_elements(22)); -- 
    cr_261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(22), ack => RPIPE_Concat_input_pipe_89_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_89_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_89_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_89_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_93_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_93_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_93_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_101_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_101_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_101_Sample/rr
      -- 
    ca_262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_89_inst_ack_1, ack => concat_CP_34_elements(23)); -- 
    rr_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(23), ack => RPIPE_Concat_input_pipe_101_inst_req_0); -- 
    rr_270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(23), ack => type_cast_93_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_93_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_93_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_93_Sample/ra
      -- 
    ra_271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_93_inst_ack_0, ack => concat_CP_34_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	74 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_93_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_93_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_93_Update/ca
      -- 
    ca_276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_93_inst_ack_1, ack => concat_CP_34_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_101_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_101_update_start_
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_101_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_101_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_101_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_101_Update/cr
      -- 
    ra_285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_101_inst_ack_0, ack => concat_CP_34_elements(26)); -- 
    cr_289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(26), ack => RPIPE_Concat_input_pipe_101_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (9) 
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_101_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_101_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_101_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_105_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_105_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_105_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_114_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_114_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_114_Sample/rr
      -- 
    ca_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_101_inst_ack_1, ack => concat_CP_34_elements(27)); -- 
    rr_298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(27), ack => type_cast_105_inst_req_0); -- 
    rr_312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(27), ack => RPIPE_Concat_input_pipe_114_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_105_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_105_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_105_Sample/ra
      -- 
    ra_299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_105_inst_ack_0, ack => concat_CP_34_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	83 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_105_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_105_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_105_Update/ca
      -- 
    ca_304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_105_inst_ack_1, ack => concat_CP_34_elements(29)); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_114_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_114_update_start_
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_114_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_114_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_114_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_114_Update/cr
      -- 
    ra_313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_114_inst_ack_0, ack => concat_CP_34_elements(30)); -- 
    cr_317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(30), ack => RPIPE_Concat_input_pipe_114_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_114_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_114_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_114_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_118_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_118_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_118_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_126_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_126_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_126_Sample/rr
      -- 
    ca_318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_114_inst_ack_1, ack => concat_CP_34_elements(31)); -- 
    rr_340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(31), ack => RPIPE_Concat_input_pipe_126_inst_req_0); -- 
    rr_326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(31), ack => type_cast_118_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_118_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_118_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_118_Sample/ra
      -- 
    ra_327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_118_inst_ack_0, ack => concat_CP_34_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	83 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_118_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_118_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_118_Update/ca
      -- 
    ca_332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_118_inst_ack_1, ack => concat_CP_34_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_126_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_126_update_start_
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_126_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_126_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_126_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_126_Update/cr
      -- 
    ra_341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_126_inst_ack_0, ack => concat_CP_34_elements(34)); -- 
    cr_345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(34), ack => RPIPE_Concat_input_pipe_126_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_126_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_126_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_126_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_130_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_130_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_130_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_139_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_139_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_139_Sample/rr
      -- 
    ca_346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_126_inst_ack_1, ack => concat_CP_34_elements(35)); -- 
    rr_354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(35), ack => type_cast_130_inst_req_0); -- 
    rr_368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(35), ack => RPIPE_Concat_input_pipe_139_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_130_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_130_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_130_Sample/ra
      -- 
    ra_355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_130_inst_ack_0, ack => concat_CP_34_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	80 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_130_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_130_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_130_Update/ca
      -- 
    ca_360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_130_inst_ack_1, ack => concat_CP_34_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_139_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_139_update_start_
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_139_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_139_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_139_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_139_Update/cr
      -- 
    ra_369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_139_inst_ack_0, ack => concat_CP_34_elements(38)); -- 
    cr_373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(38), ack => RPIPE_Concat_input_pipe_139_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_143_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_143_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_143_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_139_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_139_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_139_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_151_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_151_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_151_Sample/rr
      -- 
    ca_374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_139_inst_ack_1, ack => concat_CP_34_elements(39)); -- 
    rr_382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(39), ack => type_cast_143_inst_req_0); -- 
    rr_396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(39), ack => RPIPE_Concat_input_pipe_151_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_143_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_143_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_143_Sample/ra
      -- 
    ra_383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_143_inst_ack_0, ack => concat_CP_34_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	80 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_143_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_143_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_143_Update/ca
      -- 
    ca_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_143_inst_ack_1, ack => concat_CP_34_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_151_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_151_update_start_
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_151_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_151_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_151_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_151_Update/cr
      -- 
    ra_397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_151_inst_ack_0, ack => concat_CP_34_elements(42)); -- 
    cr_401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(42), ack => RPIPE_Concat_input_pipe_151_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	46 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_151_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_151_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_151_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_155_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_155_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_155_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_164_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_164_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_164_Sample/rr
      -- 
    ca_402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_151_inst_ack_1, ack => concat_CP_34_elements(43)); -- 
    rr_410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(43), ack => type_cast_155_inst_req_0); -- 
    rr_424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(43), ack => RPIPE_Concat_input_pipe_164_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_155_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_155_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_155_Sample/ra
      -- 
    ra_411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_0, ack => concat_CP_34_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	80 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_155_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_155_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_155_Update/ca
      -- 
    ca_416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_1, ack => concat_CP_34_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_164_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_164_update_start_
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_164_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_164_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_164_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_164_Update/cr
      -- 
    ra_425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_164_inst_ack_0, ack => concat_CP_34_elements(46)); -- 
    cr_429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(46), ack => RPIPE_Concat_input_pipe_164_inst_req_1); -- 
    -- CP-element group 47:  fork  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: 	50 
    -- CP-element group 47:  members (9) 
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_164_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_164_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_164_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_168_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_168_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_168_Sample/rr
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_176_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_176_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_176_Sample/rr
      -- 
    ca_430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_164_inst_ack_1, ack => concat_CP_34_elements(47)); -- 
    rr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(47), ack => RPIPE_Concat_input_pipe_176_inst_req_0); -- 
    rr_438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(47), ack => type_cast_168_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_168_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_168_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_168_Sample/ra
      -- 
    ra_439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_168_inst_ack_0, ack => concat_CP_34_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	80 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_168_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_168_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_168_Update/ca
      -- 
    ca_444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_168_inst_ack_1, ack => concat_CP_34_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	47 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (6) 
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_176_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_176_update_start_
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_176_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_176_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_176_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_176_Update/cr
      -- 
    ra_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_176_inst_ack_0, ack => concat_CP_34_elements(50)); -- 
    cr_457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(50), ack => RPIPE_Concat_input_pipe_176_inst_req_1); -- 
    -- CP-element group 51:  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: 	54 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_176_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_176_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_176_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_181_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_181_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_181_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_190_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_190_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_190_Sample/rr
      -- 
    ca_458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_176_inst_ack_1, ack => concat_CP_34_elements(51)); -- 
    rr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(51), ack => type_cast_181_inst_req_0); -- 
    rr_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(51), ack => RPIPE_Concat_input_pipe_190_inst_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_181_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_181_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_181_Sample/ra
      -- 
    ra_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_181_inst_ack_0, ack => concat_CP_34_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	0 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	86 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_181_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_181_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_181_Update/ca
      -- 
    ca_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_181_inst_ack_1, ack => concat_CP_34_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	51 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_190_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_190_update_start_
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_190_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_190_Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_190_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_190_Update/cr
      -- 
    ra_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_190_inst_ack_0, ack => concat_CP_34_elements(54)); -- 
    cr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(54), ack => RPIPE_Concat_input_pipe_190_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_190_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_190_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_190_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_194_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_194_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_194_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_202_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_202_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_202_Sample/rr
      -- 
    ca_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_190_inst_ack_1, ack => concat_CP_34_elements(55)); -- 
    rr_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(55), ack => type_cast_194_inst_req_0); -- 
    rr_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(55), ack => RPIPE_Concat_input_pipe_202_inst_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_194_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_194_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_194_Sample/ra
      -- 
    ra_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_0, ack => concat_CP_34_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	86 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_194_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_194_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_194_Update/ca
      -- 
    ca_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_1, ack => concat_CP_34_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	55 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_202_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_202_update_start_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_202_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_202_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_202_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_202_Update/cr
      -- 
    ra_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_202_inst_ack_0, ack => concat_CP_34_elements(58)); -- 
    cr_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(58), ack => RPIPE_Concat_input_pipe_202_inst_req_1); -- 
    -- CP-element group 59:  fork  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	62 
    -- CP-element group 59:  members (9) 
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_202_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_202_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_202_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_206_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_206_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_206_Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_215_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_215_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_215_Sample/rr
      -- 
    ca_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_202_inst_ack_1, ack => concat_CP_34_elements(59)); -- 
    rr_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(59), ack => type_cast_206_inst_req_0); -- 
    rr_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(59), ack => RPIPE_Concat_input_pipe_215_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_206_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_206_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_206_Sample/ra
      -- 
    ra_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_206_inst_ack_0, ack => concat_CP_34_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	0 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	86 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_206_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_206_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_206_Update/ca
      -- 
    ca_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_206_inst_ack_1, ack => concat_CP_34_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_215_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_215_update_start_
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_215_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_215_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_215_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_215_Update/cr
      -- 
    ra_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_215_inst_ack_0, ack => concat_CP_34_elements(62)); -- 
    cr_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(62), ack => RPIPE_Concat_input_pipe_215_inst_req_1); -- 
    -- CP-element group 63:  fork  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_215_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_215_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_215_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_219_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_219_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_219_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_227_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_227_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_227_Sample/rr
      -- 
    ca_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_215_inst_ack_1, ack => concat_CP_34_elements(63)); -- 
    rr_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(63), ack => type_cast_219_inst_req_0); -- 
    rr_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(63), ack => RPIPE_Concat_input_pipe_227_inst_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_219_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_219_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_219_Sample/ra
      -- 
    ra_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_0, ack => concat_CP_34_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	86 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_219_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_219_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_219_Update/ca
      -- 
    ca_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_1, ack => concat_CP_34_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_227_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_227_update_start_
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_227_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_227_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_227_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_227_Update/cr
      -- 
    ra_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_227_inst_ack_0, ack => concat_CP_34_elements(66)); -- 
    cr_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(66), ack => RPIPE_Concat_input_pipe_227_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: 	70 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_227_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_227_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_227_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_231_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_231_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_231_Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_240_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_240_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_240_Sample/rr
      -- 
    ca_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_227_inst_ack_1, ack => concat_CP_34_elements(67)); -- 
    rr_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(67), ack => type_cast_231_inst_req_0); -- 
    rr_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(67), ack => RPIPE_Concat_input_pipe_240_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_231_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_231_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_231_Sample/ra
      -- 
    ra_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_231_inst_ack_0, ack => concat_CP_34_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	86 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_231_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_231_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_231_Update/ca
      -- 
    ca_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_231_inst_ack_1, ack => concat_CP_34_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	67 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_240_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_240_update_start_
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_240_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_240_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_240_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_240_Update/cr
      -- 
    ra_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_240_inst_ack_0, ack => concat_CP_34_elements(70)); -- 
    cr_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(70), ack => RPIPE_Concat_input_pipe_240_inst_req_1); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_240_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_240_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/RPIPE_Concat_input_pipe_240_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_244_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_244_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_244_Sample/rr
      -- 
    ca_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_240_inst_ack_1, ack => concat_CP_34_elements(71)); -- 
    rr_606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(71), ack => type_cast_244_inst_req_0); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_244_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_244_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_244_Sample/ra
      -- 
    ra_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_244_inst_ack_0, ack => concat_CP_34_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	86 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_244_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_244_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_244_Update/ca
      -- 
    ca_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_244_inst_ack_1, ack => concat_CP_34_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	25 
    -- CP-element group 74: 	21 
    -- CP-element group 74: 	13 
    -- CP-element group 74: 	17 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_258_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_258_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_258_Sample/rr
      -- 
    rr_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(74), ack => type_cast_258_inst_req_0); -- 
    concat_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 26) := "concat_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(25) & concat_CP_34_elements(21) & concat_CP_34_elements(13) & concat_CP_34_elements(17);
      gj_concat_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_258_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_258_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_258_Sample/ra
      -- 
    ra_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_258_inst_ack_0, ack => concat_CP_34_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	0 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	86 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_258_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_258_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_258_Update/ca
      -- 
    ca_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_258_inst_ack_1, ack => concat_CP_34_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	5 
    -- CP-element group 77: 	9 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_262_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_262_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_262_Sample/rr
      -- 
    rr_634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(77), ack => type_cast_262_inst_req_0); -- 
    concat_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "concat_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(5) & concat_CP_34_elements(9);
      gj_concat_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_262_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_262_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_262_Sample/ra
      -- 
    ra_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_262_inst_ack_0, ack => concat_CP_34_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	0 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	86 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_262_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_262_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_262_Update/ca
      -- 
    ca_640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_262_inst_ack_1, ack => concat_CP_34_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	49 
    -- CP-element group 80: 	41 
    -- CP-element group 80: 	45 
    -- CP-element group 80: 	37 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_276_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_276_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_276_Sample/rr
      -- 
    rr_648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(80), ack => type_cast_276_inst_req_0); -- 
    concat_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 26) := "concat_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(49) & concat_CP_34_elements(41) & concat_CP_34_elements(45) & concat_CP_34_elements(37);
      gj_concat_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_276_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_276_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_276_Sample/ra
      -- 
    ra_649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_276_inst_ack_0, ack => concat_CP_34_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	0 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	86 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_276_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_276_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_276_Update/ca
      -- 
    ca_654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_276_inst_ack_1, ack => concat_CP_34_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	29 
    -- CP-element group 83: 	33 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_280_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_280_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_280_Sample/rr
      -- 
    rr_662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(83), ack => type_cast_280_inst_req_0); -- 
    concat_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "concat_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(29) & concat_CP_34_elements(33);
      gj_concat_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_280_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_280_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_280_Sample/ra
      -- 
    ra_663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_280_inst_ack_0, ack => concat_CP_34_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_280_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_280_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/type_cast_280_Update/ca
      -- 
    ca_668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_280_inst_ack_1, ack => concat_CP_34_elements(85)); -- 
    -- CP-element group 86:  branch  join  transition  place  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: 	82 
    -- CP-element group 86: 	53 
    -- CP-element group 86: 	57 
    -- CP-element group 86: 	61 
    -- CP-element group 86: 	65 
    -- CP-element group 86: 	69 
    -- CP-element group 86: 	73 
    -- CP-element group 86: 	76 
    -- CP-element group 86: 	79 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (10) 
      -- CP-element group 86: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314__exit__
      -- CP-element group 86: 	 branch_block_stmt_23/if_stmt_315__entry__
      -- CP-element group 86: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_314/$exit
      -- CP-element group 86: 	 branch_block_stmt_23/if_stmt_315_dead_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_23/if_stmt_315_eval_test/$entry
      -- CP-element group 86: 	 branch_block_stmt_23/if_stmt_315_eval_test/$exit
      -- CP-element group 86: 	 branch_block_stmt_23/if_stmt_315_eval_test/branch_req
      -- CP-element group 86: 	 branch_block_stmt_23/R_cmp467_316_place
      -- CP-element group 86: 	 branch_block_stmt_23/if_stmt_315_if_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_23/if_stmt_315_else_link/$entry
      -- 
    branch_req_676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(86), ack => if_stmt_315_branch_req_0); -- 
    concat_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 26) := "concat_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= concat_CP_34_elements(85) & concat_CP_34_elements(82) & concat_CP_34_elements(53) & concat_CP_34_elements(57) & concat_CP_34_elements(61) & concat_CP_34_elements(65) & concat_CP_34_elements(69) & concat_CP_34_elements(73) & concat_CP_34_elements(76) & concat_CP_34_elements(79);
      gj_concat_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	91 
    -- CP-element group 87: 	92 
    -- CP-element group 87:  members (18) 
      -- CP-element group 87: 	 branch_block_stmt_23/merge_stmt_336__exit__
      -- CP-element group 87: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371__entry__
      -- CP-element group 87: 	 branch_block_stmt_23/if_stmt_315_if_link/$exit
      -- CP-element group 87: 	 branch_block_stmt_23/if_stmt_315_if_link/if_choice_transition
      -- CP-element group 87: 	 branch_block_stmt_23/entry_bbx_xnph469
      -- CP-element group 87: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/$entry
      -- CP-element group 87: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/type_cast_357_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/type_cast_357_update_start_
      -- CP-element group 87: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/type_cast_357_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/type_cast_357_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/type_cast_357_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/type_cast_357_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_23/merge_stmt_336_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_23/entry_bbx_xnph469_PhiReq/$entry
      -- CP-element group 87: 	 branch_block_stmt_23/merge_stmt_336_PhiAck/dummy
      -- CP-element group 87: 	 branch_block_stmt_23/merge_stmt_336_PhiAck/$exit
      -- CP-element group 87: 	 branch_block_stmt_23/merge_stmt_336_PhiAck/$entry
      -- CP-element group 87: 	 branch_block_stmt_23/entry_bbx_xnph469_PhiReq/$exit
      -- 
    if_choice_transition_681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_315_branch_ack_1, ack => concat_CP_34_elements(87)); -- 
    rr_720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(87), ack => type_cast_357_inst_req_0); -- 
    cr_725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(87), ack => type_cast_357_inst_req_1); -- 
    -- CP-element group 88:  transition  place  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	439 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_23/if_stmt_315_else_link/$exit
      -- CP-element group 88: 	 branch_block_stmt_23/if_stmt_315_else_link/else_choice_transition
      -- CP-element group 88: 	 branch_block_stmt_23/entry_forx_xcond171x_xpreheader
      -- CP-element group 88: 	 branch_block_stmt_23/entry_forx_xcond171x_xpreheader_PhiReq/$entry
      -- CP-element group 88: 	 branch_block_stmt_23/entry_forx_xcond171x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_315_branch_ack_0, ack => concat_CP_34_elements(88)); -- 
    -- CP-element group 89:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	439 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	135 
    -- CP-element group 89: 	136 
    -- CP-element group 89:  members (18) 
      -- CP-element group 89: 	 branch_block_stmt_23/merge_stmt_543__exit__
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578__entry__
      -- CP-element group 89: 	 branch_block_stmt_23/if_stmt_330_if_link/$exit
      -- CP-element group 89: 	 branch_block_stmt_23/if_stmt_330_if_link/if_choice_transition
      -- CP-element group 89: 	 branch_block_stmt_23/forx_xcond171x_xpreheader_bbx_xnph465
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/$entry
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/type_cast_564_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/type_cast_564_update_start_
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/type_cast_564_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/type_cast_564_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/type_cast_564_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/type_cast_564_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_23/merge_stmt_543_PhiReqMerge
      -- CP-element group 89: 	 branch_block_stmt_23/merge_stmt_543_PhiAck/dummy
      -- CP-element group 89: 	 branch_block_stmt_23/merge_stmt_543_PhiAck/$exit
      -- CP-element group 89: 	 branch_block_stmt_23/merge_stmt_543_PhiAck/$entry
      -- CP-element group 89: 	 branch_block_stmt_23/forx_xcond171x_xpreheader_bbx_xnph465_PhiReq/$exit
      -- CP-element group 89: 	 branch_block_stmt_23/forx_xcond171x_xpreheader_bbx_xnph465_PhiReq/$entry
      -- 
    if_choice_transition_703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_330_branch_ack_1, ack => concat_CP_34_elements(89)); -- 
    rr_1079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(89), ack => type_cast_564_inst_req_0); -- 
    cr_1084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(89), ack => type_cast_564_inst_req_1); -- 
    -- CP-element group 90:  transition  place  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	439 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	452 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_23/if_stmt_330_else_link/$exit
      -- CP-element group 90: 	 branch_block_stmt_23/if_stmt_330_else_link/else_choice_transition
      -- CP-element group 90: 	 branch_block_stmt_23/forx_xcond171x_xpreheader_forx_xend231
      -- CP-element group 90: 	 branch_block_stmt_23/forx_xcond171x_xpreheader_forx_xend231_PhiReq/$exit
      -- CP-element group 90: 	 branch_block_stmt_23/forx_xcond171x_xpreheader_forx_xend231_PhiReq/$entry
      -- 
    else_choice_transition_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_330_branch_ack_0, ack => concat_CP_34_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	87 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/type_cast_357_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/type_cast_357_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/type_cast_357_Sample/ra
      -- 
    ra_721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_0, ack => concat_CP_34_elements(91)); -- 
    -- CP-element group 92:  transition  place  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	87 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	440 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371__exit__
      -- CP-element group 92: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody
      -- CP-element group 92: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/$entry
      -- CP-element group 92: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/$exit
      -- CP-element group 92: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/type_cast_357_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/type_cast_357_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_23/assign_stmt_342_to_assign_stmt_371/type_cast_357_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_374/$entry
      -- CP-element group 92: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/$entry
      -- 
    ca_726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_1, ack => concat_CP_34_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	445 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	132 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_final_index_sum_regn_Sample/ack
      -- CP-element group 93: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_final_index_sum_regn_sample_complete
      -- CP-element group 93: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_final_index_sum_regn_Sample/$exit
      -- 
    ack_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_386_index_offset_ack_0, ack => concat_CP_34_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	445 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (11) 
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_final_index_sum_regn_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_final_index_sum_regn_Update/ack
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_base_plus_offset/$entry
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_base_plus_offset/$exit
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_base_plus_offset/sum_rename_req
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_base_plus_offset/sum_rename_ack
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/addr_of_387_request/$entry
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/addr_of_387_request/req
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/addr_of_387_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_root_address_calculated
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_offset_calculated
      -- 
    ack_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_386_index_offset_ack_1, ack => concat_CP_34_elements(94)); -- 
    req_769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(94), ack => addr_of_387_final_reg_req_0); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/addr_of_387_request/$exit
      -- CP-element group 95: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/addr_of_387_request/ack
      -- CP-element group 95: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/addr_of_387_sample_completed_
      -- 
    ack_770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_387_final_reg_ack_0, ack => concat_CP_34_elements(95)); -- 
    -- CP-element group 96:  fork  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	445 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	129 
    -- CP-element group 96:  members (19) 
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/addr_of_387_complete/$exit
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/addr_of_387_complete/ack
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/addr_of_387_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_base_address_calculated
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_word_address_calculated
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_root_address_calculated
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_base_address_resized
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_base_addr_resize/$entry
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_base_addr_resize/$exit
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_base_addr_resize/base_resize_req
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_base_addr_resize/base_resize_ack
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_base_plus_offset/$entry
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_base_plus_offset/$exit
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_base_plus_offset/sum_rename_req
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_base_plus_offset/sum_rename_ack
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_word_addrgen/$entry
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_word_addrgen/$exit
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_word_addrgen/root_register_req
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_word_addrgen/root_register_ack
      -- 
    ack_775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_387_final_reg_ack_1, ack => concat_CP_34_elements(96)); -- 
    -- CP-element group 97:  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	445 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (6) 
      -- CP-element group 97: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_390_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_390_update_start_
      -- CP-element group 97: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_390_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_390_Sample/ra
      -- CP-element group 97: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_390_Update/$entry
      -- CP-element group 97: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_390_Update/cr
      -- 
    ra_784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_390_inst_ack_0, ack => concat_CP_34_elements(97)); -- 
    cr_788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(97), ack => RPIPE_Concat_input_pipe_390_inst_req_1); -- 
    -- CP-element group 98:  fork  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98: 	101 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_390_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_390_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_390_Update/ca
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_394_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_394_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_394_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_403_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_403_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_403_Sample/rr
      -- 
    ca_789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_390_inst_ack_1, ack => concat_CP_34_elements(98)); -- 
    rr_811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(98), ack => RPIPE_Concat_input_pipe_403_inst_req_0); -- 
    rr_797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(98), ack => type_cast_394_inst_req_0); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_394_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_394_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_394_Sample/ra
      -- 
    ra_798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_394_inst_ack_0, ack => concat_CP_34_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	445 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	129 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_394_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_394_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_394_Update/ca
      -- 
    ca_803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_394_inst_ack_1, ack => concat_CP_34_elements(100)); -- 
    -- CP-element group 101:  transition  input  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	98 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (6) 
      -- CP-element group 101: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_403_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_403_update_start_
      -- CP-element group 101: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_403_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_403_Sample/ra
      -- CP-element group 101: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_403_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_403_Update/cr
      -- 
    ra_812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_403_inst_ack_0, ack => concat_CP_34_elements(101)); -- 
    cr_816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(101), ack => RPIPE_Concat_input_pipe_403_inst_req_1); -- 
    -- CP-element group 102:  fork  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102: 	105 
    -- CP-element group 102:  members (9) 
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_403_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_403_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_403_Update/ca
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_407_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_407_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_407_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_421_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_421_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_421_Sample/rr
      -- 
    ca_817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_403_inst_ack_1, ack => concat_CP_34_elements(102)); -- 
    rr_839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(102), ack => RPIPE_Concat_input_pipe_421_inst_req_0); -- 
    rr_825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(102), ack => type_cast_407_inst_req_0); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_407_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_407_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_407_Sample/ra
      -- 
    ra_826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_407_inst_ack_0, ack => concat_CP_34_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	445 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	129 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_407_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_407_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_407_Update/ca
      -- 
    ca_831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_407_inst_ack_1, ack => concat_CP_34_elements(104)); -- 
    -- CP-element group 105:  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	102 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (6) 
      -- CP-element group 105: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_421_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_421_update_start_
      -- CP-element group 105: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_421_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_421_Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_421_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_421_Update/cr
      -- 
    ra_840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_421_inst_ack_0, ack => concat_CP_34_elements(105)); -- 
    cr_844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(105), ack => RPIPE_Concat_input_pipe_421_inst_req_1); -- 
    -- CP-element group 106:  fork  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106: 	109 
    -- CP-element group 106:  members (9) 
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_421_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_421_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_421_Update/ca
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_425_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_425_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_425_Sample/rr
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_439_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_439_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_439_Sample/rr
      -- 
    ca_845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_421_inst_ack_1, ack => concat_CP_34_elements(106)); -- 
    rr_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(106), ack => type_cast_425_inst_req_0); -- 
    rr_867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(106), ack => RPIPE_Concat_input_pipe_439_inst_req_0); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_425_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_425_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_425_Sample/ra
      -- 
    ra_854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_425_inst_ack_0, ack => concat_CP_34_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	445 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	129 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_425_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_425_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_425_Update/ca
      -- 
    ca_859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_425_inst_ack_1, ack => concat_CP_34_elements(108)); -- 
    -- CP-element group 109:  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	106 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (6) 
      -- CP-element group 109: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_439_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_439_update_start_
      -- CP-element group 109: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_439_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_439_Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_439_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_439_Update/cr
      -- 
    ra_868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_439_inst_ack_0, ack => concat_CP_34_elements(109)); -- 
    cr_872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(109), ack => RPIPE_Concat_input_pipe_439_inst_req_1); -- 
    -- CP-element group 110:  fork  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (9) 
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_439_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_439_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_439_Update/ca
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_443_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_443_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_443_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_457_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_457_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_457_Sample/rr
      -- 
    ca_873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_439_inst_ack_1, ack => concat_CP_34_elements(110)); -- 
    rr_881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(110), ack => type_cast_443_inst_req_0); -- 
    rr_895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(110), ack => RPIPE_Concat_input_pipe_457_inst_req_0); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_443_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_443_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_443_Sample/ra
      -- 
    ra_882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_443_inst_ack_0, ack => concat_CP_34_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	445 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	129 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_443_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_443_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_443_Update/ca
      -- 
    ca_887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_443_inst_ack_1, ack => concat_CP_34_elements(112)); -- 
    -- CP-element group 113:  transition  input  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	110 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (6) 
      -- CP-element group 113: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_457_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_457_update_start_
      -- CP-element group 113: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_457_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_457_Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_457_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_457_Update/cr
      -- 
    ra_896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_457_inst_ack_0, ack => concat_CP_34_elements(113)); -- 
    cr_900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(113), ack => RPIPE_Concat_input_pipe_457_inst_req_1); -- 
    -- CP-element group 114:  fork  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114: 	117 
    -- CP-element group 114:  members (9) 
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_457_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_457_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_457_Update/ca
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_461_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_461_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_461_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_475_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_475_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_475_Sample/rr
      -- 
    ca_901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_457_inst_ack_1, ack => concat_CP_34_elements(114)); -- 
    rr_909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(114), ack => type_cast_461_inst_req_0); -- 
    rr_923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(114), ack => RPIPE_Concat_input_pipe_475_inst_req_0); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_461_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_461_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_461_Sample/ra
      -- 
    ra_910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_461_inst_ack_0, ack => concat_CP_34_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	445 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	129 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_461_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_461_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_461_Update/ca
      -- 
    ca_915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_461_inst_ack_1, ack => concat_CP_34_elements(116)); -- 
    -- CP-element group 117:  transition  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	114 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (6) 
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_475_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_475_update_start_
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_475_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_475_Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_475_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_475_Update/cr
      -- 
    ra_924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_475_inst_ack_0, ack => concat_CP_34_elements(117)); -- 
    cr_928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(117), ack => RPIPE_Concat_input_pipe_475_inst_req_1); -- 
    -- CP-element group 118:  fork  transition  input  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	121 
    -- CP-element group 118:  members (9) 
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_475_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_475_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_475_Update/ca
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_479_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_479_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_479_Sample/rr
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_493_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_493_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_493_Sample/rr
      -- 
    ca_929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_475_inst_ack_1, ack => concat_CP_34_elements(118)); -- 
    rr_937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(118), ack => type_cast_479_inst_req_0); -- 
    rr_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(118), ack => RPIPE_Concat_input_pipe_493_inst_req_0); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_479_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_479_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_479_Sample/ra
      -- 
    ra_938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_479_inst_ack_0, ack => concat_CP_34_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	445 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	129 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_479_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_479_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_479_Update/ca
      -- 
    ca_943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_479_inst_ack_1, ack => concat_CP_34_elements(120)); -- 
    -- CP-element group 121:  transition  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	118 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (6) 
      -- CP-element group 121: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_493_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_493_update_start_
      -- CP-element group 121: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_493_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_493_Sample/ra
      -- CP-element group 121: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_493_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_493_Update/cr
      -- 
    ra_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_493_inst_ack_0, ack => concat_CP_34_elements(121)); -- 
    cr_956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(121), ack => RPIPE_Concat_input_pipe_493_inst_req_1); -- 
    -- CP-element group 122:  fork  transition  input  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122: 	125 
    -- CP-element group 122:  members (9) 
      -- CP-element group 122: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_493_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_493_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_493_Update/ca
      -- CP-element group 122: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_497_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_497_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_497_Sample/rr
      -- CP-element group 122: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_511_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_511_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_511_Sample/rr
      -- 
    ca_957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_493_inst_ack_1, ack => concat_CP_34_elements(122)); -- 
    rr_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(122), ack => type_cast_497_inst_req_0); -- 
    rr_979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(122), ack => RPIPE_Concat_input_pipe_511_inst_req_0); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_497_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_497_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_497_Sample/ra
      -- 
    ra_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_497_inst_ack_0, ack => concat_CP_34_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	445 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	129 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_497_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_497_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_497_Update/ca
      -- 
    ca_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_497_inst_ack_1, ack => concat_CP_34_elements(124)); -- 
    -- CP-element group 125:  transition  input  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	122 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (6) 
      -- CP-element group 125: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_511_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_511_update_start_
      -- CP-element group 125: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_511_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_511_Sample/ra
      -- CP-element group 125: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_511_Update/$entry
      -- CP-element group 125: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_511_Update/cr
      -- 
    ra_980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_511_inst_ack_0, ack => concat_CP_34_elements(125)); -- 
    cr_984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(125), ack => RPIPE_Concat_input_pipe_511_inst_req_1); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (6) 
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_511_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_511_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_511_Update/ca
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_515_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_515_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_515_Sample/rr
      -- 
    ca_985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_511_inst_ack_1, ack => concat_CP_34_elements(126)); -- 
    rr_993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(126), ack => type_cast_515_inst_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_515_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_515_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_515_Sample/ra
      -- 
    ra_994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_515_inst_ack_0, ack => concat_CP_34_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	445 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_515_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_515_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_515_Update/ca
      -- 
    ca_999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_515_inst_ack_1, ack => concat_CP_34_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	104 
    -- CP-element group 129: 	108 
    -- CP-element group 129: 	112 
    -- CP-element group 129: 	116 
    -- CP-element group 129: 	120 
    -- CP-element group 129: 	124 
    -- CP-element group 129: 	128 
    -- CP-element group 129: 	100 
    -- CP-element group 129: 	96 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (9) 
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Sample/ptr_deref_523_Split/$entry
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Sample/ptr_deref_523_Split/$exit
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Sample/ptr_deref_523_Split/split_req
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Sample/ptr_deref_523_Split/split_ack
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Sample/word_access_start/$entry
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Sample/word_access_start/word_0/$entry
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Sample/word_access_start/word_0/rr
      -- 
    rr_1037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(129), ack => ptr_deref_523_store_0_req_0); -- 
    concat_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= concat_CP_34_elements(104) & concat_CP_34_elements(108) & concat_CP_34_elements(112) & concat_CP_34_elements(116) & concat_CP_34_elements(120) & concat_CP_34_elements(124) & concat_CP_34_elements(128) & concat_CP_34_elements(100) & concat_CP_34_elements(96);
      gj_concat_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (5) 
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Sample/word_access_start/$exit
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Sample/word_access_start/word_0/$exit
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Sample/word_access_start/word_0/ra
      -- 
    ra_1038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_523_store_0_ack_0, ack => concat_CP_34_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	445 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (5) 
      -- CP-element group 131: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Update/word_access_complete/$exit
      -- CP-element group 131: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Update/word_access_complete/word_0/$exit
      -- CP-element group 131: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Update/word_access_complete/word_0/ca
      -- 
    ca_1049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_523_store_0_ack_1, ack => concat_CP_34_elements(131)); -- 
    -- CP-element group 132:  branch  join  transition  place  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: 	93 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (10) 
      -- CP-element group 132: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536__exit__
      -- CP-element group 132: 	 branch_block_stmt_23/if_stmt_537__entry__
      -- CP-element group 132: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/$exit
      -- CP-element group 132: 	 branch_block_stmt_23/if_stmt_537_dead_link/$entry
      -- CP-element group 132: 	 branch_block_stmt_23/if_stmt_537_eval_test/$entry
      -- CP-element group 132: 	 branch_block_stmt_23/if_stmt_537_eval_test/$exit
      -- CP-element group 132: 	 branch_block_stmt_23/if_stmt_537_eval_test/branch_req
      -- CP-element group 132: 	 branch_block_stmt_23/R_exitcond2_538_place
      -- CP-element group 132: 	 branch_block_stmt_23/if_stmt_537_if_link/$entry
      -- CP-element group 132: 	 branch_block_stmt_23/if_stmt_537_else_link/$entry
      -- 
    branch_req_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(132), ack => if_stmt_537_branch_req_0); -- 
    concat_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(131) & concat_CP_34_elements(93);
      gj_concat_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  merge  transition  place  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	439 
    -- CP-element group 133:  members (13) 
      -- CP-element group 133: 	 branch_block_stmt_23/merge_stmt_321__exit__
      -- CP-element group 133: 	 branch_block_stmt_23/forx_xcond171x_xpreheaderx_xloopexit_forx_xcond171x_xpreheader
      -- CP-element group 133: 	 branch_block_stmt_23/if_stmt_537_if_link/$exit
      -- CP-element group 133: 	 branch_block_stmt_23/if_stmt_537_if_link/if_choice_transition
      -- CP-element group 133: 	 branch_block_stmt_23/forx_xbody_forx_xcond171x_xpreheaderx_xloopexit
      -- CP-element group 133: 	 branch_block_stmt_23/forx_xbody_forx_xcond171x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 133: 	 branch_block_stmt_23/forx_xbody_forx_xcond171x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 133: 	 branch_block_stmt_23/merge_stmt_321_PhiReqMerge
      -- CP-element group 133: 	 branch_block_stmt_23/merge_stmt_321_PhiAck/$entry
      -- CP-element group 133: 	 branch_block_stmt_23/merge_stmt_321_PhiAck/$exit
      -- CP-element group 133: 	 branch_block_stmt_23/merge_stmt_321_PhiAck/dummy
      -- CP-element group 133: 	 branch_block_stmt_23/forx_xcond171x_xpreheaderx_xloopexit_forx_xcond171x_xpreheader_PhiReq/$entry
      -- CP-element group 133: 	 branch_block_stmt_23/forx_xcond171x_xpreheaderx_xloopexit_forx_xcond171x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_537_branch_ack_1, ack => concat_CP_34_elements(133)); -- 
    -- CP-element group 134:  fork  transition  place  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	441 
    -- CP-element group 134: 	442 
    -- CP-element group 134:  members (12) 
      -- CP-element group 134: 	 branch_block_stmt_23/if_stmt_537_else_link/$exit
      -- CP-element group 134: 	 branch_block_stmt_23/if_stmt_537_else_link/else_choice_transition
      -- CP-element group 134: 	 branch_block_stmt_23/forx_xbody_forx_xbody
      -- CP-element group 134: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/type_cast_380/SplitProtocol/Update/cr
      -- CP-element group 134: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 134: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/$entry
      -- CP-element group 134: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/type_cast_380/SplitProtocol/Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/type_cast_380/SplitProtocol/Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/type_cast_380/SplitProtocol/Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/type_cast_380/SplitProtocol/$entry
      -- CP-element group 134: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/type_cast_380/$entry
      -- CP-element group 134: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/$entry
      -- 
    else_choice_transition_1066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_537_branch_ack_0, ack => concat_CP_34_elements(134)); -- 
    cr_2759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(134), ack => type_cast_380_inst_req_1); -- 
    rr_2754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(134), ack => type_cast_380_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	89 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/type_cast_564_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/type_cast_564_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/type_cast_564_Sample/ra
      -- 
    ra_1080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_564_inst_ack_0, ack => concat_CP_34_elements(135)); -- 
    -- CP-element group 136:  transition  place  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	89 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	446 
    -- CP-element group 136:  members (9) 
      -- CP-element group 136: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578__exit__
      -- CP-element group 136: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177
      -- CP-element group 136: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/$exit
      -- CP-element group 136: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/type_cast_564_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/type_cast_564_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_23/assign_stmt_549_to_assign_stmt_578/type_cast_564_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/$entry
      -- CP-element group 136: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_581/$entry
      -- CP-element group 136: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/$entry
      -- 
    ca_1085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_564_inst_ack_1, ack => concat_CP_34_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	451 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	176 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_final_index_sum_regn_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_final_index_sum_regn_Sample/ack
      -- CP-element group 137: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_final_index_sum_regn_sample_complete
      -- 
    ack_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_593_index_offset_ack_0, ack => concat_CP_34_elements(137)); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	451 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (11) 
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_base_plus_offset/sum_rename_ack
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_base_plus_offset/sum_rename_req
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_base_plus_offset/$exit
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_base_plus_offset/$entry
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_final_index_sum_regn_Update/ack
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_final_index_sum_regn_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/addr_of_594_request/req
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/addr_of_594_request/$entry
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/addr_of_594_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_root_address_calculated
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_offset_calculated
      -- 
    ack_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_593_index_offset_ack_1, ack => concat_CP_34_elements(138)); -- 
    req_1128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(138), ack => addr_of_594_final_reg_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/addr_of_594_request/ack
      -- CP-element group 139: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/addr_of_594_request/$exit
      -- CP-element group 139: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/addr_of_594_sample_completed_
      -- 
    ack_1129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_594_final_reg_ack_0, ack => concat_CP_34_elements(139)); -- 
    -- CP-element group 140:  fork  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	451 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	173 
    -- CP-element group 140:  members (19) 
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_base_plus_offset/$exit
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_base_plus_offset/$entry
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_base_address_resized
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_base_addr_resize/base_resize_ack
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_base_addr_resize/base_resize_req
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_base_addr_resize/$exit
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_base_addr_resize/$entry
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_root_address_calculated
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_word_address_calculated
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_base_address_calculated
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_word_addrgen/root_register_ack
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_word_addrgen/root_register_req
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_word_addrgen/$exit
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_word_addrgen/$entry
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_base_plus_offset/sum_rename_ack
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_base_plus_offset/sum_rename_req
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/addr_of_594_complete/ack
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/addr_of_594_complete/$exit
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/addr_of_594_update_completed_
      -- 
    ack_1134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_594_final_reg_ack_1, ack => concat_CP_34_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	451 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_597_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_597_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_597_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_597_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_597_update_start_
      -- CP-element group 141: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_597_sample_completed_
      -- 
    ra_1143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_597_inst_ack_0, ack => concat_CP_34_elements(141)); -- 
    cr_1147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(141), ack => RPIPE_Concat_input_pipe_597_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_610_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_610_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_610_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_601_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_601_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_601_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_597_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_597_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_597_update_completed_
      -- 
    ca_1148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_597_inst_ack_1, ack => concat_CP_34_elements(142)); -- 
    rr_1156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(142), ack => type_cast_601_inst_req_0); -- 
    rr_1170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(142), ack => RPIPE_Concat_input_pipe_610_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_601_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_601_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_601_sample_completed_
      -- 
    ra_1157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_601_inst_ack_0, ack => concat_CP_34_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	451 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	173 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_601_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_601_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_601_update_completed_
      -- 
    ca_1162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_601_inst_ack_1, ack => concat_CP_34_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_610_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_610_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_610_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_610_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_610_update_start_
      -- CP-element group 145: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_610_sample_completed_
      -- 
    ra_1171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_610_inst_ack_0, ack => concat_CP_34_elements(145)); -- 
    cr_1175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(145), ack => RPIPE_Concat_input_pipe_610_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_628_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_610_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_610_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_614_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_614_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_614_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_610_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_628_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_628_Sample/$entry
      -- 
    ca_1176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_610_inst_ack_1, ack => concat_CP_34_elements(146)); -- 
    rr_1184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(146), ack => type_cast_614_inst_req_0); -- 
    rr_1198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(146), ack => RPIPE_Concat_input_pipe_628_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_614_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_614_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_614_Sample/$exit
      -- 
    ra_1185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_614_inst_ack_0, ack => concat_CP_34_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	451 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	173 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_614_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_614_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_614_update_completed_
      -- 
    ca_1190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_614_inst_ack_1, ack => concat_CP_34_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_628_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_628_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_628_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_628_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_628_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_628_update_start_
      -- 
    ra_1199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_628_inst_ack_0, ack => concat_CP_34_elements(149)); -- 
    cr_1203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(149), ack => RPIPE_Concat_input_pipe_628_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_646_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_646_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_646_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_632_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_632_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_632_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_628_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_628_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_628_update_completed_
      -- 
    ca_1204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_628_inst_ack_1, ack => concat_CP_34_elements(150)); -- 
    rr_1212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(150), ack => type_cast_632_inst_req_0); -- 
    rr_1226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(150), ack => RPIPE_Concat_input_pipe_646_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_632_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_632_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_632_sample_completed_
      -- 
    ra_1213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_632_inst_ack_0, ack => concat_CP_34_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	451 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	173 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_632_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_632_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_632_update_completed_
      -- 
    ca_1218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_632_inst_ack_1, ack => concat_CP_34_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_646_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_646_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_646_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_646_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_646_update_start_
      -- CP-element group 153: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_646_sample_completed_
      -- 
    ra_1227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_646_inst_ack_0, ack => concat_CP_34_elements(153)); -- 
    cr_1231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(153), ack => RPIPE_Concat_input_pipe_646_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_646_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_646_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_646_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_664_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_664_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_664_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_650_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_650_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_650_sample_start_
      -- 
    ca_1232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_646_inst_ack_1, ack => concat_CP_34_elements(154)); -- 
    rr_1240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(154), ack => type_cast_650_inst_req_0); -- 
    rr_1254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(154), ack => RPIPE_Concat_input_pipe_664_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_650_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_650_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_650_sample_completed_
      -- 
    ra_1241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_650_inst_ack_0, ack => concat_CP_34_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	451 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	173 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_650_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_650_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_650_update_completed_
      -- 
    ca_1246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_650_inst_ack_1, ack => concat_CP_34_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_664_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_664_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_664_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_664_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_664_update_start_
      -- CP-element group 157: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_664_sample_completed_
      -- 
    ra_1255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_664_inst_ack_0, ack => concat_CP_34_elements(157)); -- 
    cr_1259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(157), ack => RPIPE_Concat_input_pipe_664_inst_req_1); -- 
    -- CP-element group 158:  fork  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	161 
    -- CP-element group 158:  members (9) 
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_668_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_668_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_668_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_664_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_664_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_664_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_682_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_682_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_682_sample_start_
      -- 
    ca_1260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_664_inst_ack_1, ack => concat_CP_34_elements(158)); -- 
    rr_1282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(158), ack => RPIPE_Concat_input_pipe_682_inst_req_0); -- 
    rr_1268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(158), ack => type_cast_668_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_668_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_668_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_668_sample_completed_
      -- 
    ra_1269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_668_inst_ack_0, ack => concat_CP_34_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	451 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	173 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_668_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_668_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_668_update_completed_
      -- 
    ca_1274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_668_inst_ack_1, ack => concat_CP_34_elements(160)); -- 
    -- CP-element group 161:  transition  input  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	158 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (6) 
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_682_Update/cr
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_682_Update/$entry
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_682_Sample/ra
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_682_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_682_update_start_
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_682_sample_completed_
      -- 
    ra_1283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_682_inst_ack_0, ack => concat_CP_34_elements(161)); -- 
    cr_1287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(161), ack => RPIPE_Concat_input_pipe_682_inst_req_1); -- 
    -- CP-element group 162:  fork  transition  input  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162: 	165 
    -- CP-element group 162:  members (9) 
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_686_Sample/rr
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_686_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_686_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_700_Sample/rr
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_700_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_682_Update/ca
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_682_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_700_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_682_update_completed_
      -- 
    ca_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_682_inst_ack_1, ack => concat_CP_34_elements(162)); -- 
    rr_1296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(162), ack => type_cast_686_inst_req_0); -- 
    rr_1310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(162), ack => RPIPE_Concat_input_pipe_700_inst_req_0); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_686_Sample/ra
      -- CP-element group 163: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_686_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_686_sample_completed_
      -- 
    ra_1297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_686_inst_ack_0, ack => concat_CP_34_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	451 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	173 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_686_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_686_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_686_Update/ca
      -- 
    ca_1302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_686_inst_ack_1, ack => concat_CP_34_elements(164)); -- 
    -- CP-element group 165:  transition  input  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	162 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (6) 
      -- CP-element group 165: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_700_Update/cr
      -- CP-element group 165: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_700_Update/$entry
      -- CP-element group 165: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_700_Sample/ra
      -- CP-element group 165: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_700_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_700_update_start_
      -- CP-element group 165: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_700_sample_completed_
      -- 
    ra_1311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_700_inst_ack_0, ack => concat_CP_34_elements(165)); -- 
    cr_1315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(165), ack => RPIPE_Concat_input_pipe_700_inst_req_1); -- 
    -- CP-element group 166:  fork  transition  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166: 	169 
    -- CP-element group 166:  members (9) 
      -- CP-element group 166: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_704_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_718_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_700_Update/ca
      -- CP-element group 166: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_700_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_718_Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_700_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_718_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_704_Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_704_Sample/$entry
      -- 
    ca_1316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_700_inst_ack_1, ack => concat_CP_34_elements(166)); -- 
    rr_1324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(166), ack => type_cast_704_inst_req_0); -- 
    rr_1338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(166), ack => RPIPE_Concat_input_pipe_718_inst_req_0); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_704_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_704_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_704_Sample/$exit
      -- 
    ra_1325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_704_inst_ack_0, ack => concat_CP_34_elements(167)); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	451 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	173 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_704_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_704_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_704_Update/$exit
      -- 
    ca_1330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_704_inst_ack_1, ack => concat_CP_34_elements(168)); -- 
    -- CP-element group 169:  transition  input  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	166 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (6) 
      -- CP-element group 169: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_718_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_718_Update/cr
      -- CP-element group 169: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_718_Update/$entry
      -- CP-element group 169: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_718_Sample/ra
      -- CP-element group 169: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_718_update_start_
      -- CP-element group 169: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_718_sample_completed_
      -- 
    ra_1339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_718_inst_ack_0, ack => concat_CP_34_elements(169)); -- 
    cr_1343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(169), ack => RPIPE_Concat_input_pipe_718_inst_req_1); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (6) 
      -- CP-element group 170: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_722_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_718_Update/ca
      -- CP-element group 170: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_718_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_718_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_722_Sample/rr
      -- CP-element group 170: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_722_Sample/$entry
      -- 
    ca_1344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_718_inst_ack_1, ack => concat_CP_34_elements(170)); -- 
    rr_1352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(170), ack => type_cast_722_inst_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_722_Sample/ra
      -- CP-element group 171: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_722_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_722_sample_completed_
      -- 
    ra_1353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_722_inst_ack_0, ack => concat_CP_34_elements(171)); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	451 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_722_Update/ca
      -- CP-element group 172: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_722_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_722_update_completed_
      -- 
    ca_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_722_inst_ack_1, ack => concat_CP_34_elements(172)); -- 
    -- CP-element group 173:  join  transition  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	160 
    -- CP-element group 173: 	172 
    -- CP-element group 173: 	168 
    -- CP-element group 173: 	140 
    -- CP-element group 173: 	144 
    -- CP-element group 173: 	148 
    -- CP-element group 173: 	152 
    -- CP-element group 173: 	156 
    -- CP-element group 173: 	164 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (9) 
      -- CP-element group 173: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Sample/ptr_deref_730_Split/split_ack
      -- CP-element group 173: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Sample/ptr_deref_730_Split/split_req
      -- CP-element group 173: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Sample/ptr_deref_730_Split/$exit
      -- CP-element group 173: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Sample/ptr_deref_730_Split/$entry
      -- CP-element group 173: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Sample/word_access_start/word_0/rr
      -- CP-element group 173: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Sample/word_access_start/word_0/$entry
      -- CP-element group 173: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Sample/word_access_start/$entry
      -- 
    rr_1396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(173), ack => ptr_deref_730_store_0_req_0); -- 
    concat_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= concat_CP_34_elements(160) & concat_CP_34_elements(172) & concat_CP_34_elements(168) & concat_CP_34_elements(140) & concat_CP_34_elements(144) & concat_CP_34_elements(148) & concat_CP_34_elements(152) & concat_CP_34_elements(156) & concat_CP_34_elements(164);
      gj_concat_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (5) 
      -- CP-element group 174: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Sample/word_access_start/word_0/ra
      -- CP-element group 174: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Sample/word_access_start/word_0/$exit
      -- CP-element group 174: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Sample/word_access_start/$exit
      -- 
    ra_1397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_730_store_0_ack_0, ack => concat_CP_34_elements(174)); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	451 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (5) 
      -- CP-element group 175: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Update/word_access_complete/word_0/ca
      -- CP-element group 175: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Update/word_access_complete/word_0/$exit
      -- CP-element group 175: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Update/word_access_complete/$exit
      -- CP-element group 175: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Update/$exit
      -- 
    ca_1408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_730_store_0_ack_1, ack => concat_CP_34_elements(175)); -- 
    -- CP-element group 176:  branch  join  transition  place  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: 	137 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (10) 
      -- CP-element group 176: 	 branch_block_stmt_23/if_stmt_744_eval_test/branch_req
      -- CP-element group 176: 	 branch_block_stmt_23/if_stmt_744_eval_test/$exit
      -- CP-element group 176: 	 branch_block_stmt_23/if_stmt_744_eval_test/$entry
      -- CP-element group 176: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743__exit__
      -- CP-element group 176: 	 branch_block_stmt_23/if_stmt_744__entry__
      -- CP-element group 176: 	 branch_block_stmt_23/if_stmt_744_dead_link/$entry
      -- CP-element group 176: 	 branch_block_stmt_23/if_stmt_744_else_link/$entry
      -- CP-element group 176: 	 branch_block_stmt_23/if_stmt_744_if_link/$entry
      -- CP-element group 176: 	 branch_block_stmt_23/R_exitcond_745_place
      -- CP-element group 176: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/$exit
      -- 
    branch_req_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(176), ack => if_stmt_744_branch_req_0); -- 
    concat_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(175) & concat_CP_34_elements(137);
      gj_concat_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  merge  transition  place  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	452 
    -- CP-element group 177:  members (13) 
      -- CP-element group 177: 	 branch_block_stmt_23/merge_stmt_750__exit__
      -- CP-element group 177: 	 branch_block_stmt_23/forx_xend231x_xloopexit_forx_xend231
      -- CP-element group 177: 	 branch_block_stmt_23/forx_xbody177_forx_xend231x_xloopexit
      -- CP-element group 177: 	 branch_block_stmt_23/merge_stmt_750_PhiAck/$exit
      -- CP-element group 177: 	 branch_block_stmt_23/if_stmt_744_if_link/if_choice_transition
      -- CP-element group 177: 	 branch_block_stmt_23/if_stmt_744_if_link/$exit
      -- CP-element group 177: 	 branch_block_stmt_23/merge_stmt_750_PhiReqMerge
      -- CP-element group 177: 	 branch_block_stmt_23/forx_xbody177_forx_xend231x_xloopexit_PhiReq/$entry
      -- CP-element group 177: 	 branch_block_stmt_23/forx_xbody177_forx_xend231x_xloopexit_PhiReq/$exit
      -- CP-element group 177: 	 branch_block_stmt_23/merge_stmt_750_PhiAck/$entry
      -- CP-element group 177: 	 branch_block_stmt_23/forx_xend231x_xloopexit_forx_xend231_PhiReq/$exit
      -- CP-element group 177: 	 branch_block_stmt_23/forx_xend231x_xloopexit_forx_xend231_PhiReq/$entry
      -- CP-element group 177: 	 branch_block_stmt_23/merge_stmt_750_PhiAck/dummy
      -- 
    if_choice_transition_1421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_744_branch_ack_1, ack => concat_CP_34_elements(177)); -- 
    -- CP-element group 178:  fork  transition  place  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	447 
    -- CP-element group 178: 	448 
    -- CP-element group 178:  members (12) 
      -- CP-element group 178: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/$entry
      -- CP-element group 178: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177
      -- CP-element group 178: 	 branch_block_stmt_23/if_stmt_744_else_link/else_choice_transition
      -- CP-element group 178: 	 branch_block_stmt_23/if_stmt_744_else_link/$exit
      -- CP-element group 178: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/$entry
      -- CP-element group 178: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/$entry
      -- CP-element group 178: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/type_cast_587/$entry
      -- CP-element group 178: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/type_cast_587/SplitProtocol/$entry
      -- CP-element group 178: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/type_cast_587/SplitProtocol/Update/cr
      -- CP-element group 178: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/type_cast_587/SplitProtocol/Update/$entry
      -- CP-element group 178: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/type_cast_587/SplitProtocol/Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/type_cast_587/SplitProtocol/Sample/$entry
      -- 
    else_choice_transition_1425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_744_branch_ack_0, ack => concat_CP_34_elements(178)); -- 
    cr_2813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(178), ack => type_cast_587_inst_req_1); -- 
    rr_2808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(178), ack => type_cast_587_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	452 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_23/call_stmt_755/call_stmt_755_Sample/cra
      -- CP-element group 179: 	 branch_block_stmt_23/call_stmt_755/call_stmt_755_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_23/call_stmt_755/call_stmt_755_sample_completed_
      -- 
    cra_1439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_755_call_ack_0, ack => concat_CP_34_elements(179)); -- 
    -- CP-element group 180:  transition  place  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	452 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (10) 
      -- CP-element group 180: 	 branch_block_stmt_23/call_stmt_755/call_stmt_755_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_23/assign_stmt_762_to_assign_stmt_783/$exit
      -- CP-element group 180: 	 branch_block_stmt_23/call_stmt_755__exit__
      -- CP-element group 180: 	 branch_block_stmt_23/assign_stmt_762_to_assign_stmt_783__entry__
      -- CP-element group 180: 	 branch_block_stmt_23/assign_stmt_762_to_assign_stmt_783__exit__
      -- CP-element group 180: 	 branch_block_stmt_23/do_while_stmt_784__entry__
      -- CP-element group 180: 	 branch_block_stmt_23/assign_stmt_762_to_assign_stmt_783/$entry
      -- CP-element group 180: 	 branch_block_stmt_23/call_stmt_755/call_stmt_755_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_23/call_stmt_755/$exit
      -- CP-element group 180: 	 branch_block_stmt_23/call_stmt_755/call_stmt_755_Update/cca
      -- 
    cca_1444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_755_call_ack_1, ack => concat_CP_34_elements(180)); -- 
    -- CP-element group 181:  transition  place  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	187 
    -- CP-element group 181:  members (2) 
      -- CP-element group 181: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784__entry__
      -- CP-element group 181: 	 branch_block_stmt_23/do_while_stmt_784/$entry
      -- 
    concat_CP_34_elements(181) <= concat_CP_34_elements(180);
    -- CP-element group 182:  merge  place  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	333 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784__exit__
      -- 
    -- Element group concat_CP_34_elements(182) is bound as output of CP function.
    -- CP-element group 183:  merge  place  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	186 
    -- CP-element group 183:  members (1) 
      -- CP-element group 183: 	 branch_block_stmt_23/do_while_stmt_784/loop_back
      -- 
    -- Element group concat_CP_34_elements(183) is bound as output of CP function.
    -- CP-element group 184:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	189 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	331 
    -- CP-element group 184: 	332 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_23/do_while_stmt_784/condition_done
      -- CP-element group 184: 	 branch_block_stmt_23/do_while_stmt_784/loop_exit/$entry
      -- CP-element group 184: 	 branch_block_stmt_23/do_while_stmt_784/loop_taken/$entry
      -- 
    concat_CP_34_elements(184) <= concat_CP_34_elements(189);
    -- CP-element group 185:  branch  place  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	330 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_23/do_while_stmt_784/loop_body_done
      -- 
    concat_CP_34_elements(185) <= concat_CP_34_elements(330);
    -- CP-element group 186:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	183 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	198 
    -- CP-element group 186: 	217 
    -- CP-element group 186: 	236 
    -- CP-element group 186: 	255 
    -- CP-element group 186:  members (1) 
      -- CP-element group 186: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/back_edge_to_loop_body
      -- 
    concat_CP_34_elements(186) <= concat_CP_34_elements(183);
    -- CP-element group 187:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	181 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	200 
    -- CP-element group 187: 	219 
    -- CP-element group 187: 	238 
    -- CP-element group 187: 	257 
    -- CP-element group 187:  members (1) 
      -- CP-element group 187: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/first_time_through_loop_body
      -- 
    concat_CP_34_elements(187) <= concat_CP_34_elements(181);
    -- CP-element group 188:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	194 
    -- CP-element group 188: 	195 
    -- CP-element group 188: 	211 
    -- CP-element group 188: 	212 
    -- CP-element group 188: 	230 
    -- CP-element group 188: 	231 
    -- CP-element group 188: 	321 
    -- CP-element group 188: 	325 
    -- CP-element group 188: 	329 
    -- CP-element group 188: 	249 
    -- CP-element group 188: 	250 
    -- CP-element group 188: 	269 
    -- CP-element group 188: 	270 
    -- CP-element group 188: 	284 
    -- CP-element group 188: 	285 
    -- CP-element group 188: 	299 
    -- CP-element group 188: 	300 
    -- CP-element group 188:  members (2) 
      -- CP-element group 188: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/loop_body_start
      -- CP-element group 188: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/$entry
      -- 
    -- Element group concat_CP_34_elements(188) is bound as output of CP function.
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	193 
    -- CP-element group 189: 	197 
    -- CP-element group 189: 	324 
    -- CP-element group 189: 	328 
    -- CP-element group 189: 	329 
    -- CP-element group 189: 	254 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	184 
    -- CP-element group 189:  members (1) 
      -- CP-element group 189: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/condition_evaluated
      -- 
    condition_evaluated_1462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(189), ack => do_while_stmt_784_branch_req_0); -- 
    concat_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(193) & concat_CP_34_elements(197) & concat_CP_34_elements(324) & concat_CP_34_elements(328) & concat_CP_34_elements(329) & concat_CP_34_elements(254);
      gj_concat_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	194 
    -- CP-element group 190: 	211 
    -- CP-element group 190: 	230 
    -- CP-element group 190: 	249 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	193 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	213 
    -- CP-element group 190: 	232 
    -- CP-element group 190: 	251 
    -- CP-element group 190:  members (2) 
      -- CP-element group 190: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_sample_start__ps
      -- CP-element group 190: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/aggregated_phi_sample_req
      -- 
    concat_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(194) & concat_CP_34_elements(211) & concat_CP_34_elements(230) & concat_CP_34_elements(249) & concat_CP_34_elements(193);
      gj_concat_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	196 
    -- CP-element group 191: 	214 
    -- CP-element group 191: 	233 
    -- CP-element group 191: 	252 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	322 
    -- CP-element group 191: 	330 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	194 
    -- CP-element group 191: 	211 
    -- CP-element group 191: 	230 
    -- CP-element group 191: 	249 
    -- CP-element group 191:  members (5) 
      -- CP-element group 191: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/aggregated_phi_sample_ack
      -- CP-element group 191: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_sample_completed_
      -- 
    concat_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(196) & concat_CP_34_elements(214) & concat_CP_34_elements(233) & concat_CP_34_elements(252);
      gj_concat_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	195 
    -- CP-element group 192: 	212 
    -- CP-element group 192: 	231 
    -- CP-element group 192: 	250 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	215 
    -- CP-element group 192: 	234 
    -- CP-element group 192: 	253 
    -- CP-element group 192:  members (2) 
      -- CP-element group 192: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_update_start__ps
      -- CP-element group 192: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/aggregated_phi_update_req
      -- 
    concat_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(195) & concat_CP_34_elements(212) & concat_CP_34_elements(231) & concat_CP_34_elements(250);
      gj_concat_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	197 
    -- CP-element group 193: 	216 
    -- CP-element group 193: 	235 
    -- CP-element group 193: 	254 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	189 
    -- CP-element group 193: marked-successors 
    -- CP-element group 193: 	190 
    -- CP-element group 193:  members (1) 
      -- CP-element group 193: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/aggregated_phi_update_ack
      -- 
    concat_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(197) & concat_CP_34_elements(216) & concat_CP_34_elements(235) & concat_CP_34_elements(254);
      gj_concat_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  join  transition  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	188 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	191 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	190 
    -- CP-element group 194:  members (1) 
      -- CP-element group 194: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_sample_start_
      -- 
    concat_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(191);
      gj_concat_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  join  transition  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	188 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	197 
    -- CP-element group 195: 	301 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	192 
    -- CP-element group 195:  members (1) 
      -- CP-element group 195: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_update_start_
      -- 
    concat_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(197) & concat_CP_34_elements(301);
      gj_concat_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  join  transition  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	191 
    -- CP-element group 196:  members (1) 
      -- CP-element group 196: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(196) is bound as output of CP function.
    -- CP-element group 197:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	189 
    -- CP-element group 197: 	193 
    -- CP-element group 197: 	301 
    -- CP-element group 197: marked-successors 
    -- CP-element group 197: 	195 
    -- CP-element group 197:  members (15) 
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_index_computed_1
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_index_resize_1/index_resize_ack
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_index_scale_1/$entry
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_index_resize_1/$entry
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_final_index_sum_regn_Sample/req
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_index_scale_1/scale_rename_req
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_index_resize_1/$exit
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_index_scale_1/scale_rename_ack
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_index_resize_1/index_resize_req
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_final_index_sum_regn_Sample/$entry
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_index_scale_1/$exit
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_update_completed__ps
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_index_scaled_1
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_index_resized_1
      -- 
    req_1888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(197), ack => array_obj_ref_845_index_offset_req_0); -- 
    -- Element group concat_CP_34_elements(197) is bound as output of CP function.
    -- CP-element group 198:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	186 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_loopback_trigger
      -- 
    concat_CP_34_elements(198) <= concat_CP_34_elements(186);
    -- CP-element group 199:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (2) 
      -- CP-element group 199: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_loopback_sample_req
      -- CP-element group 199: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_loopback_sample_req_ps
      -- 
    phi_stmt_786_loopback_sample_req_1477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_786_loopback_sample_req_1477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(199), ack => phi_stmt_786_req_1); -- 
    -- Element group concat_CP_34_elements(199) is bound as output of CP function.
    -- CP-element group 200:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	187 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_entry_trigger
      -- 
    concat_CP_34_elements(200) <= concat_CP_34_elements(187);
    -- CP-element group 201:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (2) 
      -- CP-element group 201: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_entry_sample_req
      -- CP-element group 201: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_entry_sample_req_ps
      -- 
    phi_stmt_786_entry_sample_req_1480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_786_entry_sample_req_1480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(201), ack => phi_stmt_786_req_0); -- 
    -- Element group concat_CP_34_elements(201) is bound as output of CP function.
    -- CP-element group 202:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (2) 
      -- CP-element group 202: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_phi_mux_ack
      -- CP-element group 202: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_786_phi_mux_ack_ps
      -- 
    phi_stmt_786_phi_mux_ack_1483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_786_ack_0, ack => concat_CP_34_elements(202)); -- 
    -- CP-element group 203:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (4) 
      -- CP-element group 203: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_out_init_788_sample_start__ps
      -- CP-element group 203: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_out_init_788_sample_completed__ps
      -- CP-element group 203: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_out_init_788_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_out_init_788_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(203) is bound as output of CP function.
    -- CP-element group 204:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (2) 
      -- CP-element group 204: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_out_init_788_update_start__ps
      -- CP-element group 204: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_out_init_788_update_start_
      -- 
    -- Element group concat_CP_34_elements(204) is bound as output of CP function.
    -- CP-element group 205:  join  transition  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	206 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (1) 
      -- CP-element group 205: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_out_init_788_update_completed__ps
      -- 
    concat_CP_34_elements(205) <= concat_CP_34_elements(206);
    -- CP-element group 206:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	205 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_out_init_788_update_completed_
      -- 
    -- Element group concat_CP_34_elements(206) is a control-delay.
    cp_element_206_delay: control_delay_element  generic map(name => " 206_delay", delay_value => 1)  port map(req => concat_CP_34_elements(204), ack => concat_CP_34_elements(206), clk => clk, reset =>reset);
    -- CP-element group 207:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (4) 
      -- CP-element group 207: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_sample_start__ps
      -- CP-element group 207: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_Sample/req
      -- 
    req_1504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(207), ack => next_add_out_899_789_buf_req_0); -- 
    -- Element group concat_CP_34_elements(207) is bound as output of CP function.
    -- CP-element group 208:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (4) 
      -- CP-element group 208: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_update_start__ps
      -- CP-element group 208: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_update_start_
      -- CP-element group 208: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_Update/req
      -- 
    req_1509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(208), ack => next_add_out_899_789_buf_req_1); -- 
    -- Element group concat_CP_34_elements(208) is bound as output of CP function.
    -- CP-element group 209:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (4) 
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_sample_completed__ps
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_sample_completed_
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_Sample/ack
      -- 
    ack_1505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_out_899_789_buf_ack_0, ack => concat_CP_34_elements(209)); -- 
    -- CP-element group 210:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (4) 
      -- CP-element group 210: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_update_completed__ps
      -- CP-element group 210: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_out_789_Update/ack
      -- 
    ack_1510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_out_899_789_buf_ack_1, ack => concat_CP_34_elements(210)); -- 
    -- CP-element group 211:  join  transition  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	188 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	191 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	190 
    -- CP-element group 211:  members (1) 
      -- CP-element group 211: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_sample_start_
      -- 
    concat_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(191);
      gj_concat_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  join  transition  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	188 
    -- CP-element group 212: marked-predecessors 
    -- CP-element group 212: 	216 
    -- CP-element group 212: 	271 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	192 
    -- CP-element group 212:  members (1) 
      -- CP-element group 212: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_update_start_
      -- 
    concat_cp_element_group_212: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_212"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(216) & concat_CP_34_elements(271);
      gj_concat_cp_element_group_212 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 213:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	190 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (1) 
      -- CP-element group 213: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_sample_start__ps
      -- 
    concat_CP_34_elements(213) <= concat_CP_34_elements(190);
    -- CP-element group 214:  join  transition  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	191 
    -- CP-element group 214:  members (1) 
      -- CP-element group 214: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(214) is bound as output of CP function.
    -- CP-element group 215:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	192 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (1) 
      -- CP-element group 215: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_update_start__ps
      -- 
    concat_CP_34_elements(215) <= concat_CP_34_elements(192);
    -- CP-element group 216:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	193 
    -- CP-element group 216: 	271 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	212 
    -- CP-element group 216:  members (15) 
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_update_completed__ps
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_index_resized_1
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_index_scaled_1
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_index_computed_1
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_index_resize_1/$entry
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_index_resize_1/$exit
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_index_resize_1/index_resize_req
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_index_resize_1/index_resize_ack
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_index_scale_1/$entry
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_index_scale_1/$exit
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_index_scale_1/scale_rename_req
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_index_scale_1/scale_rename_ack
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_final_index_sum_regn_Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_final_index_sum_regn_Sample/req
      -- 
    req_1668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(216), ack => array_obj_ref_813_index_offset_req_0); -- 
    -- Element group concat_CP_34_elements(216) is bound as output of CP function.
    -- CP-element group 217:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	186 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (1) 
      -- CP-element group 217: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_loopback_trigger
      -- 
    concat_CP_34_elements(217) <= concat_CP_34_elements(186);
    -- CP-element group 218:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: successors 
    -- CP-element group 218:  members (2) 
      -- CP-element group 218: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_loopback_sample_req
      -- CP-element group 218: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_loopback_sample_req_ps
      -- 
    phi_stmt_790_loopback_sample_req_1521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_790_loopback_sample_req_1521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(218), ack => phi_stmt_790_req_1); -- 
    -- Element group concat_CP_34_elements(218) is bound as output of CP function.
    -- CP-element group 219:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	187 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (1) 
      -- CP-element group 219: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_entry_trigger
      -- 
    concat_CP_34_elements(219) <= concat_CP_34_elements(187);
    -- CP-element group 220:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (2) 
      -- CP-element group 220: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_entry_sample_req
      -- CP-element group 220: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_entry_sample_req_ps
      -- 
    phi_stmt_790_entry_sample_req_1524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_790_entry_sample_req_1524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(220), ack => phi_stmt_790_req_0); -- 
    -- Element group concat_CP_34_elements(220) is bound as output of CP function.
    -- CP-element group 221:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (2) 
      -- CP-element group 221: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_phi_mux_ack
      -- CP-element group 221: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_790_phi_mux_ack_ps
      -- 
    phi_stmt_790_phi_mux_ack_1527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_790_ack_0, ack => concat_CP_34_elements(221)); -- 
    -- CP-element group 222:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: successors 
    -- CP-element group 222:  members (4) 
      -- CP-element group 222: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp1_init_792_sample_start__ps
      -- CP-element group 222: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp1_init_792_sample_completed__ps
      -- CP-element group 222: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp1_init_792_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp1_init_792_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(222) is bound as output of CP function.
    -- CP-element group 223:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (2) 
      -- CP-element group 223: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp1_init_792_update_start__ps
      -- CP-element group 223: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp1_init_792_update_start_
      -- 
    -- Element group concat_CP_34_elements(223) is bound as output of CP function.
    -- CP-element group 224:  join  transition  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	225 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (1) 
      -- CP-element group 224: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp1_init_792_update_completed__ps
      -- 
    concat_CP_34_elements(224) <= concat_CP_34_elements(225);
    -- CP-element group 225:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	224 
    -- CP-element group 225:  members (1) 
      -- CP-element group 225: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp1_init_792_update_completed_
      -- 
    -- Element group concat_CP_34_elements(225) is a control-delay.
    cp_element_225_delay: control_delay_element  generic map(name => " 225_delay", delay_value => 1)  port map(req => concat_CP_34_elements(223), ack => concat_CP_34_elements(225), clk => clk, reset =>reset);
    -- CP-element group 226:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (4) 
      -- CP-element group 226: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_sample_start__ps
      -- CP-element group 226: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_Sample/req
      -- 
    req_1548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(226), ack => next_add_inp1_886_793_buf_req_0); -- 
    -- Element group concat_CP_34_elements(226) is bound as output of CP function.
    -- CP-element group 227:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (4) 
      -- CP-element group 227: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_update_start__ps
      -- CP-element group 227: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_update_start_
      -- CP-element group 227: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_Update/req
      -- 
    req_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(227), ack => next_add_inp1_886_793_buf_req_1); -- 
    -- Element group concat_CP_34_elements(227) is bound as output of CP function.
    -- CP-element group 228:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (4) 
      -- CP-element group 228: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_sample_completed__ps
      -- CP-element group 228: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_Sample/ack
      -- 
    ack_1549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_inp1_886_793_buf_ack_0, ack => concat_CP_34_elements(228)); -- 
    -- CP-element group 229:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229:  members (4) 
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_update_completed__ps
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp1_793_Update/ack
      -- 
    ack_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_inp1_886_793_buf_ack_1, ack => concat_CP_34_elements(229)); -- 
    -- CP-element group 230:  join  transition  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	188 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	191 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	190 
    -- CP-element group 230:  members (1) 
      -- CP-element group 230: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_sample_start_
      -- 
    concat_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(191);
      gj_concat_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  join  transition  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	188 
    -- CP-element group 231: marked-predecessors 
    -- CP-element group 231: 	235 
    -- CP-element group 231: 	286 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	192 
    -- CP-element group 231:  members (1) 
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_update_start_
      -- 
    concat_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(235) & concat_CP_34_elements(286);
      gj_concat_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	190 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (1) 
      -- CP-element group 232: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_sample_start__ps
      -- 
    concat_CP_34_elements(232) <= concat_CP_34_elements(190);
    -- CP-element group 233:  join  transition  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	191 
    -- CP-element group 233:  members (1) 
      -- CP-element group 233: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(233) is bound as output of CP function.
    -- CP-element group 234:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	192 
    -- CP-element group 234: successors 
    -- CP-element group 234:  members (1) 
      -- CP-element group 234: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_update_start__ps
      -- 
    concat_CP_34_elements(234) <= concat_CP_34_elements(192);
    -- CP-element group 235:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	193 
    -- CP-element group 235: 	286 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	231 
    -- CP-element group 235:  members (15) 
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_update_completed_
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_update_completed__ps
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_index_resized_1
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_index_scaled_1
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_index_computed_1
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_index_resize_1/$entry
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_index_resize_1/$exit
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_index_resize_1/index_resize_req
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_index_resize_1/index_resize_ack
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_index_scale_1/$entry
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_index_scale_1/$exit
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_index_scale_1/scale_rename_req
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_index_scale_1/scale_rename_ack
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_final_index_sum_regn_Sample/$entry
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_final_index_sum_regn_Sample/req
      -- 
    req_1778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(235), ack => array_obj_ref_829_index_offset_req_0); -- 
    -- Element group concat_CP_34_elements(235) is bound as output of CP function.
    -- CP-element group 236:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	186 
    -- CP-element group 236: successors 
    -- CP-element group 236:  members (1) 
      -- CP-element group 236: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_loopback_trigger
      -- 
    concat_CP_34_elements(236) <= concat_CP_34_elements(186);
    -- CP-element group 237:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (2) 
      -- CP-element group 237: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_loopback_sample_req
      -- CP-element group 237: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_loopback_sample_req_ps
      -- 
    phi_stmt_794_loopback_sample_req_1565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_794_loopback_sample_req_1565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(237), ack => phi_stmt_794_req_1); -- 
    -- Element group concat_CP_34_elements(237) is bound as output of CP function.
    -- CP-element group 238:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	187 
    -- CP-element group 238: successors 
    -- CP-element group 238:  members (1) 
      -- CP-element group 238: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_entry_trigger
      -- 
    concat_CP_34_elements(238) <= concat_CP_34_elements(187);
    -- CP-element group 239:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (2) 
      -- CP-element group 239: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_entry_sample_req
      -- CP-element group 239: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_entry_sample_req_ps
      -- 
    phi_stmt_794_entry_sample_req_1568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_794_entry_sample_req_1568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(239), ack => phi_stmt_794_req_0); -- 
    -- Element group concat_CP_34_elements(239) is bound as output of CP function.
    -- CP-element group 240:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (2) 
      -- CP-element group 240: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_phi_mux_ack
      -- CP-element group 240: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_794_phi_mux_ack_ps
      -- 
    phi_stmt_794_phi_mux_ack_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_794_ack_0, ack => concat_CP_34_elements(240)); -- 
    -- CP-element group 241:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (4) 
      -- CP-element group 241: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp2_init_796_sample_start__ps
      -- CP-element group 241: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp2_init_796_sample_completed__ps
      -- CP-element group 241: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp2_init_796_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp2_init_796_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(241) is bound as output of CP function.
    -- CP-element group 242:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (2) 
      -- CP-element group 242: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp2_init_796_update_start__ps
      -- CP-element group 242: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp2_init_796_update_start_
      -- 
    -- Element group concat_CP_34_elements(242) is bound as output of CP function.
    -- CP-element group 243:  join  transition  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	244 
    -- CP-element group 243: successors 
    -- CP-element group 243:  members (1) 
      -- CP-element group 243: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp2_init_796_update_completed__ps
      -- 
    concat_CP_34_elements(243) <= concat_CP_34_elements(244);
    -- CP-element group 244:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	243 
    -- CP-element group 244:  members (1) 
      -- CP-element group 244: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_add_inp2_init_796_update_completed_
      -- 
    -- Element group concat_CP_34_elements(244) is a control-delay.
    cp_element_244_delay: control_delay_element  generic map(name => " 244_delay", delay_value => 1)  port map(req => concat_CP_34_elements(242), ack => concat_CP_34_elements(244), clk => clk, reset =>reset);
    -- CP-element group 245:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (4) 
      -- CP-element group 245: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_sample_start__ps
      -- CP-element group 245: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_Sample/req
      -- 
    req_1592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(245), ack => next_add_inp2_894_797_buf_req_0); -- 
    -- Element group concat_CP_34_elements(245) is bound as output of CP function.
    -- CP-element group 246:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (4) 
      -- CP-element group 246: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_update_start__ps
      -- CP-element group 246: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_update_start_
      -- CP-element group 246: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_Update/req
      -- 
    req_1597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(246), ack => next_add_inp2_894_797_buf_req_1); -- 
    -- Element group concat_CP_34_elements(246) is bound as output of CP function.
    -- CP-element group 247:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247:  members (4) 
      -- CP-element group 247: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_sample_completed__ps
      -- CP-element group 247: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_Sample/ack
      -- 
    ack_1593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_inp2_894_797_buf_ack_0, ack => concat_CP_34_elements(247)); -- 
    -- CP-element group 248:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (4) 
      -- CP-element group 248: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_update_completed__ps
      -- CP-element group 248: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_add_inp2_797_Update/ack
      -- 
    ack_1598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_inp2_894_797_buf_ack_1, ack => concat_CP_34_elements(248)); -- 
    -- CP-element group 249:  join  transition  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	188 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	191 
    -- CP-element group 249: 	324 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	190 
    -- CP-element group 249:  members (1) 
      -- CP-element group 249: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_sample_start_
      -- 
    concat_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(191) & concat_CP_34_elements(324);
      gj_concat_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  join  transition  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	188 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	311 
    -- CP-element group 250: 	254 
    -- CP-element group 250: 	277 
    -- CP-element group 250: 	292 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	192 
    -- CP-element group 250:  members (1) 
      -- CP-element group 250: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_update_start_
      -- 
    concat_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(311) & concat_CP_34_elements(254) & concat_CP_34_elements(277) & concat_CP_34_elements(292);
      gj_concat_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	190 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (1) 
      -- CP-element group 251: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_sample_start__ps
      -- 
    concat_CP_34_elements(251) <= concat_CP_34_elements(190);
    -- CP-element group 252:  join  transition  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	191 
    -- CP-element group 252:  members (1) 
      -- CP-element group 252: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(252) is bound as output of CP function.
    -- CP-element group 253:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	192 
    -- CP-element group 253: successors 
    -- CP-element group 253:  members (1) 
      -- CP-element group 253: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_update_start__ps
      -- 
    concat_CP_34_elements(253) <= concat_CP_34_elements(192);
    -- CP-element group 254:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	189 
    -- CP-element group 254: 	193 
    -- CP-element group 254: 	309 
    -- CP-element group 254: 	275 
    -- CP-element group 254: 	290 
    -- CP-element group 254: marked-successors 
    -- CP-element group 254: 	250 
    -- CP-element group 254:  members (2) 
      -- CP-element group 254: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_update_completed__ps
      -- 
    -- Element group concat_CP_34_elements(254) is bound as output of CP function.
    -- CP-element group 255:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	186 
    -- CP-element group 255: successors 
    -- CP-element group 255:  members (1) 
      -- CP-element group 255: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_loopback_trigger
      -- 
    concat_CP_34_elements(255) <= concat_CP_34_elements(186);
    -- CP-element group 256:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: successors 
    -- CP-element group 256:  members (2) 
      -- CP-element group 256: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_loopback_sample_req
      -- CP-element group 256: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_loopback_sample_req_ps
      -- 
    phi_stmt_798_loopback_sample_req_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_798_loopback_sample_req_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(256), ack => phi_stmt_798_req_1); -- 
    -- Element group concat_CP_34_elements(256) is bound as output of CP function.
    -- CP-element group 257:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	187 
    -- CP-element group 257: successors 
    -- CP-element group 257:  members (1) 
      -- CP-element group 257: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_entry_trigger
      -- 
    concat_CP_34_elements(257) <= concat_CP_34_elements(187);
    -- CP-element group 258:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: successors 
    -- CP-element group 258:  members (2) 
      -- CP-element group 258: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_entry_sample_req
      -- CP-element group 258: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_entry_sample_req_ps
      -- 
    phi_stmt_798_entry_sample_req_1612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_798_entry_sample_req_1612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(258), ack => phi_stmt_798_req_0); -- 
    -- Element group concat_CP_34_elements(258) is bound as output of CP function.
    -- CP-element group 259:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: successors 
    -- CP-element group 259:  members (2) 
      -- CP-element group 259: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_phi_mux_ack_ps
      -- CP-element group 259: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/phi_stmt_798_phi_mux_ack
      -- 
    phi_stmt_798_phi_mux_ack_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_798_ack_0, ack => concat_CP_34_elements(259)); -- 
    -- CP-element group 260:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: successors 
    -- CP-element group 260:  members (4) 
      -- CP-element group 260: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_count_inp1_init_800_sample_start__ps
      -- CP-element group 260: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_count_inp1_init_800_sample_completed__ps
      -- CP-element group 260: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_count_inp1_init_800_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_count_inp1_init_800_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(260) is bound as output of CP function.
    -- CP-element group 261:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (2) 
      -- CP-element group 261: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_count_inp1_init_800_update_start__ps
      -- CP-element group 261: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_count_inp1_init_800_update_start_
      -- 
    -- Element group concat_CP_34_elements(261) is bound as output of CP function.
    -- CP-element group 262:  join  transition  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	263 
    -- CP-element group 262: successors 
    -- CP-element group 262:  members (1) 
      -- CP-element group 262: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_count_inp1_init_800_update_completed__ps
      -- 
    concat_CP_34_elements(262) <= concat_CP_34_elements(263);
    -- CP-element group 263:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	262 
    -- CP-element group 263:  members (1) 
      -- CP-element group 263: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_count_inp1_init_800_update_completed_
      -- 
    -- Element group concat_CP_34_elements(263) is a control-delay.
    cp_element_263_delay: control_delay_element  generic map(name => " 263_delay", delay_value => 1)  port map(req => concat_CP_34_elements(261), ack => concat_CP_34_elements(263), clk => clk, reset =>reset);
    -- CP-element group 264:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (4) 
      -- CP-element group 264: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_sample_start__ps
      -- CP-element group 264: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_Sample/req
      -- 
    req_1636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(264), ack => next_count_inp1_878_801_buf_req_0); -- 
    -- Element group concat_CP_34_elements(264) is bound as output of CP function.
    -- CP-element group 265:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (4) 
      -- CP-element group 265: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_update_start__ps
      -- CP-element group 265: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_update_start_
      -- CP-element group 265: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_Update/$entry
      -- CP-element group 265: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_Update/req
      -- 
    req_1641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(265), ack => next_count_inp1_878_801_buf_req_1); -- 
    -- Element group concat_CP_34_elements(265) is bound as output of CP function.
    -- CP-element group 266:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266:  members (4) 
      -- CP-element group 266: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_sample_completed__ps
      -- CP-element group 266: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_Sample/ack
      -- 
    ack_1637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_inp1_878_801_buf_ack_0, ack => concat_CP_34_elements(266)); -- 
    -- CP-element group 267:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267:  members (4) 
      -- CP-element group 267: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_update_completed__ps
      -- CP-element group 267: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_update_completed_
      -- CP-element group 267: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/R_next_count_inp1_801_Update/ack
      -- 
    ack_1642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_inp1_878_801_buf_ack_1, ack => concat_CP_34_elements(267)); -- 
    -- CP-element group 268:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	272 
    -- CP-element group 268: marked-predecessors 
    -- CP-element group 268: 	273 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	273 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_814_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_814_request/$entry
      -- CP-element group 268: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_814_request/req
      -- 
    req_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(268), ack => addr_of_814_final_reg_req_0); -- 
    concat_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(272) & concat_CP_34_elements(273);
      gj_concat_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	188 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	274 
    -- CP-element group 269: 	281 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	274 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_814_update_start_
      -- CP-element group 269: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_814_complete/$entry
      -- CP-element group 269: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_814_complete/req
      -- 
    req_1688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(269), ack => addr_of_814_final_reg_req_1); -- 
    concat_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(274) & concat_CP_34_elements(281);
      gj_concat_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	188 
    -- CP-element group 270: marked-predecessors 
    -- CP-element group 270: 	272 
    -- CP-element group 270: 	273 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_final_index_sum_regn_update_start
      -- CP-element group 270: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_final_index_sum_regn_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_final_index_sum_regn_Update/req
      -- 
    req_1673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(270), ack => array_obj_ref_813_index_offset_req_1); -- 
    concat_cp_element_group_270: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_270"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(272) & concat_CP_34_elements(273);
      gj_concat_cp_element_group_270 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(270), clk => clk, reset => reset); --
    end block;
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	216 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	330 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	212 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_final_index_sum_regn_sample_complete
      -- CP-element group 271: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_final_index_sum_regn_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_final_index_sum_regn_Sample/ack
      -- 
    ack_1669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_813_index_offset_ack_0, ack => concat_CP_34_elements(271)); -- 
    -- CP-element group 272:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	268 
    -- CP-element group 272: marked-successors 
    -- CP-element group 272: 	270 
    -- CP-element group 272:  members (8) 
      -- CP-element group 272: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_root_address_calculated
      -- CP-element group 272: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_offset_calculated
      -- CP-element group 272: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_final_index_sum_regn_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_final_index_sum_regn_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_base_plus_offset/$entry
      -- CP-element group 272: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_base_plus_offset/$exit
      -- CP-element group 272: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_base_plus_offset/sum_rename_req
      -- CP-element group 272: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_813_base_plus_offset/sum_rename_ack
      -- 
    ack_1674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_813_index_offset_ack_1, ack => concat_CP_34_elements(272)); -- 
    -- CP-element group 273:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	268 
    -- CP-element group 273: successors 
    -- CP-element group 273: marked-successors 
    -- CP-element group 273: 	268 
    -- CP-element group 273: 	270 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_814_sample_completed_
      -- CP-element group 273: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_814_request/$exit
      -- CP-element group 273: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_814_request/ack
      -- 
    ack_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_814_final_reg_ack_0, ack => concat_CP_34_elements(273)); -- 
    -- CP-element group 274:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	269 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	279 
    -- CP-element group 274: marked-successors 
    -- CP-element group 274: 	269 
    -- CP-element group 274:  members (19) 
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_814_update_completed_
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_814_complete/$exit
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_814_complete/ack
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_base_address_calculated
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_word_address_calculated
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_root_address_calculated
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_base_address_resized
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_base_addr_resize/$entry
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_base_addr_resize/$exit
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_base_addr_resize/base_resize_req
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_base_addr_resize/base_resize_ack
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_base_plus_offset/$entry
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_base_plus_offset/$exit
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_base_plus_offset/sum_rename_req
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_base_plus_offset/sum_rename_ack
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_word_addrgen/$entry
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_word_addrgen/$exit
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_word_addrgen/root_register_req
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_word_addrgen/root_register_ack
      -- 
    ack_1689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_814_final_reg_ack_1, ack => concat_CP_34_elements(274)); -- 
    -- CP-element group 275:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	254 
    -- CP-element group 275: marked-predecessors 
    -- CP-element group 275: 	277 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	277 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_818_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_818_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_818_Sample/req
      -- 
    req_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(275), ack => W_cmp_816_delayed_6_0_816_inst_req_0); -- 
    concat_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(254) & concat_CP_34_elements(277);
      gj_concat_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: 	281 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	278 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_818_update_start_
      -- CP-element group 276: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_818_Update/$entry
      -- CP-element group 276: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_818_Update/req
      -- 
    req_1702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(276), ack => W_cmp_816_delayed_6_0_816_inst_req_1); -- 
    concat_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(278) & concat_CP_34_elements(281);
      gj_concat_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	275 
    -- CP-element group 277: successors 
    -- CP-element group 277: marked-successors 
    -- CP-element group 277: 	250 
    -- CP-element group 277: 	275 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_818_sample_completed_
      -- CP-element group 277: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_818_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_818_Sample/ack
      -- 
    ack_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_cmp_816_delayed_6_0_816_inst_ack_0, ack => concat_CP_34_elements(277)); -- 
    -- CP-element group 278:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	276 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_818_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_818_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_818_Update/ack
      -- 
    ack_1703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_cmp_816_delayed_6_0_816_inst_ack_1, ack => concat_CP_34_elements(278)); -- 
    -- CP-element group 279:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	274 
    -- CP-element group 279: 	278 
    -- CP-element group 279: marked-predecessors 
    -- CP-element group 279: 	281 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	281 
    -- CP-element group 279:  members (5) 
      -- CP-element group 279: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_sample_start_
      -- CP-element group 279: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Sample/$entry
      -- CP-element group 279: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Sample/word_access_start/$entry
      -- CP-element group 279: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Sample/word_access_start/word_0/$entry
      -- CP-element group 279: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Sample/word_access_start/word_0/rr
      -- 
    rr_1736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(279), ack => ptr_deref_822_load_0_req_0); -- 
    concat_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(274) & concat_CP_34_elements(278) & concat_CP_34_elements(281);
      gj_concat_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: marked-predecessors 
    -- CP-element group 280: 	315 
    -- CP-element group 280: 	282 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	282 
    -- CP-element group 280:  members (5) 
      -- CP-element group 280: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_update_start_
      -- CP-element group 280: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Update/$entry
      -- CP-element group 280: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Update/word_access_complete/$entry
      -- CP-element group 280: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Update/word_access_complete/word_0/$entry
      -- CP-element group 280: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Update/word_access_complete/word_0/cr
      -- 
    cr_1747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(280), ack => ptr_deref_822_load_0_req_1); -- 
    concat_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(315) & concat_CP_34_elements(282);
      gj_concat_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	279 
    -- CP-element group 281: successors 
    -- CP-element group 281: marked-successors 
    -- CP-element group 281: 	269 
    -- CP-element group 281: 	276 
    -- CP-element group 281: 	279 
    -- CP-element group 281:  members (5) 
      -- CP-element group 281: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Sample/word_access_start/$exit
      -- CP-element group 281: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Sample/word_access_start/word_0/$exit
      -- CP-element group 281: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Sample/word_access_start/word_0/ra
      -- 
    ra_1737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_822_load_0_ack_0, ack => concat_CP_34_elements(281)); -- 
    -- CP-element group 282:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	280 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	313 
    -- CP-element group 282: marked-successors 
    -- CP-element group 282: 	280 
    -- CP-element group 282:  members (9) 
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Update/word_access_complete/$exit
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Update/word_access_complete/word_0/$exit
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Update/word_access_complete/word_0/ca
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Update/ptr_deref_822_Merge/$entry
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Update/ptr_deref_822_Merge/$exit
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Update/ptr_deref_822_Merge/merge_req
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_822_Update/ptr_deref_822_Merge/merge_ack
      -- 
    ca_1748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_822_load_0_ack_1, ack => concat_CP_34_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	287 
    -- CP-element group 283: marked-predecessors 
    -- CP-element group 283: 	288 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	288 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_830_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_830_request/$entry
      -- CP-element group 283: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_830_request/req
      -- 
    req_1793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(283), ack => addr_of_830_final_reg_req_0); -- 
    concat_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(287) & concat_CP_34_elements(288);
      gj_concat_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	188 
    -- CP-element group 284: marked-predecessors 
    -- CP-element group 284: 	289 
    -- CP-element group 284: 	296 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	289 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_830_update_start_
      -- CP-element group 284: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_830_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_830_complete/req
      -- 
    req_1798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(284), ack => addr_of_830_final_reg_req_1); -- 
    concat_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(289) & concat_CP_34_elements(296);
      gj_concat_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	188 
    -- CP-element group 285: marked-predecessors 
    -- CP-element group 285: 	287 
    -- CP-element group 285: 	288 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_final_index_sum_regn_update_start
      -- CP-element group 285: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_final_index_sum_regn_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_final_index_sum_regn_Update/req
      -- 
    req_1783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(285), ack => array_obj_ref_829_index_offset_req_1); -- 
    concat_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(287) & concat_CP_34_elements(288);
      gj_concat_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	235 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	330 
    -- CP-element group 286: marked-successors 
    -- CP-element group 286: 	231 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_final_index_sum_regn_sample_complete
      -- CP-element group 286: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_final_index_sum_regn_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_final_index_sum_regn_Sample/ack
      -- 
    ack_1779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_829_index_offset_ack_0, ack => concat_CP_34_elements(286)); -- 
    -- CP-element group 287:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	283 
    -- CP-element group 287: marked-successors 
    -- CP-element group 287: 	285 
    -- CP-element group 287:  members (8) 
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_root_address_calculated
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_offset_calculated
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_final_index_sum_regn_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_final_index_sum_regn_Update/ack
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_base_plus_offset/$entry
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_base_plus_offset/$exit
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_base_plus_offset/sum_rename_req
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_829_base_plus_offset/sum_rename_ack
      -- 
    ack_1784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_829_index_offset_ack_1, ack => concat_CP_34_elements(287)); -- 
    -- CP-element group 288:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	283 
    -- CP-element group 288: successors 
    -- CP-element group 288: marked-successors 
    -- CP-element group 288: 	283 
    -- CP-element group 288: 	285 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_830_sample_completed_
      -- CP-element group 288: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_830_request/$exit
      -- CP-element group 288: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_830_request/ack
      -- 
    ack_1794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_830_final_reg_ack_0, ack => concat_CP_34_elements(288)); -- 
    -- CP-element group 289:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	284 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	294 
    -- CP-element group 289: marked-successors 
    -- CP-element group 289: 	284 
    -- CP-element group 289:  members (19) 
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_830_update_completed_
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_830_complete/$exit
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_830_complete/ack
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_base_address_calculated
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_word_address_calculated
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_root_address_calculated
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_base_address_resized
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_base_addr_resize/$entry
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_base_addr_resize/$exit
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_base_addr_resize/base_resize_req
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_base_addr_resize/base_resize_ack
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_base_plus_offset/$entry
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_base_plus_offset/$exit
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_base_plus_offset/sum_rename_req
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_base_plus_offset/sum_rename_ack
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_word_addrgen/$entry
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_word_addrgen/$exit
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_word_addrgen/root_register_req
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_word_addrgen/root_register_ack
      -- 
    ack_1799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_830_final_reg_ack_1, ack => concat_CP_34_elements(289)); -- 
    -- CP-element group 290:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	254 
    -- CP-element group 290: marked-predecessors 
    -- CP-element group 290: 	292 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_834_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_834_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_834_Sample/req
      -- 
    req_1807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(290), ack => W_cmp_829_delayed_6_0_832_inst_req_0); -- 
    concat_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(254) & concat_CP_34_elements(292);
      gj_concat_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: marked-predecessors 
    -- CP-element group 291: 	293 
    -- CP-element group 291: 	296 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_834_update_start_
      -- CP-element group 291: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_834_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_834_Update/req
      -- 
    req_1812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(291), ack => W_cmp_829_delayed_6_0_832_inst_req_1); -- 
    concat_cp_element_group_291: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_291"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(293) & concat_CP_34_elements(296);
      gj_concat_cp_element_group_291 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(291), clk => clk, reset => reset); --
    end block;
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	250 
    -- CP-element group 292: 	290 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_834_sample_completed_
      -- CP-element group 292: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_834_Sample/$exit
      -- CP-element group 292: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_834_Sample/ack
      -- 
    ack_1808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_cmp_829_delayed_6_0_832_inst_ack_0, ack => concat_CP_34_elements(292)); -- 
    -- CP-element group 293:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293: marked-successors 
    -- CP-element group 293: 	291 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_834_update_completed_
      -- CP-element group 293: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_834_Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_834_Update/ack
      -- 
    ack_1813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_cmp_829_delayed_6_0_832_inst_ack_1, ack => concat_CP_34_elements(293)); -- 
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	289 
    -- CP-element group 294: 	293 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	296 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (5) 
      -- CP-element group 294: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Sample/word_access_start/$entry
      -- CP-element group 294: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Sample/word_access_start/word_0/$entry
      -- CP-element group 294: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Sample/word_access_start/word_0/rr
      -- 
    rr_1846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(294), ack => ptr_deref_838_load_0_req_0); -- 
    concat_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(289) & concat_CP_34_elements(293) & concat_CP_34_elements(296);
      gj_concat_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: marked-predecessors 
    -- CP-element group 295: 	315 
    -- CP-element group 295: 	297 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	297 
    -- CP-element group 295:  members (5) 
      -- CP-element group 295: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_update_start_
      -- CP-element group 295: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Update/word_access_complete/$entry
      -- CP-element group 295: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Update/word_access_complete/word_0/$entry
      -- CP-element group 295: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Update/word_access_complete/word_0/cr
      -- 
    cr_1857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(295), ack => ptr_deref_838_load_0_req_1); -- 
    concat_cp_element_group_295: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_295"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(315) & concat_CP_34_elements(297);
      gj_concat_cp_element_group_295 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(295), clk => clk, reset => reset); --
    end block;
    -- CP-element group 296:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	284 
    -- CP-element group 296: 	291 
    -- CP-element group 296: 	294 
    -- CP-element group 296:  members (5) 
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_sample_completed_
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Sample/$exit
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Sample/word_access_start/$exit
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Sample/word_access_start/word_0/$exit
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Sample/word_access_start/word_0/ra
      -- 
    ra_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_838_load_0_ack_0, ack => concat_CP_34_elements(296)); -- 
    -- CP-element group 297:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	295 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	313 
    -- CP-element group 297: marked-successors 
    -- CP-element group 297: 	295 
    -- CP-element group 297:  members (9) 
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_update_completed_
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Update/$exit
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Update/word_access_complete/$exit
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Update/word_access_complete/word_0/$exit
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Update/word_access_complete/word_0/ca
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Update/ptr_deref_838_Merge/$entry
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Update/ptr_deref_838_Merge/$exit
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Update/ptr_deref_838_Merge/merge_req
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_838_Update/ptr_deref_838_Merge/merge_ack
      -- 
    ca_1858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_838_load_0_ack_1, ack => concat_CP_34_elements(297)); -- 
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	302 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	303 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	303 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_846_request/$entry
      -- CP-element group 298: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_846_request/req
      -- CP-element group 298: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_846_sample_start_
      -- 
    req_1903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(298), ack => addr_of_846_final_reg_req_0); -- 
    concat_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(302) & concat_CP_34_elements(303);
      gj_concat_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	188 
    -- CP-element group 299: marked-predecessors 
    -- CP-element group 299: 	307 
    -- CP-element group 299: 	304 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	304 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_846_complete/$entry
      -- CP-element group 299: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_846_complete/req
      -- CP-element group 299: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_846_update_start_
      -- 
    req_1908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(299), ack => addr_of_846_final_reg_req_1); -- 
    concat_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(307) & concat_CP_34_elements(304);
      gj_concat_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	188 
    -- CP-element group 300: marked-predecessors 
    -- CP-element group 300: 	302 
    -- CP-element group 300: 	303 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	302 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_final_index_sum_regn_update_start
      -- CP-element group 300: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_final_index_sum_regn_Update/$entry
      -- CP-element group 300: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_final_index_sum_regn_Update/req
      -- 
    req_1893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(300), ack => array_obj_ref_845_index_offset_req_1); -- 
    concat_cp_element_group_300: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_300"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(302) & concat_CP_34_elements(303);
      gj_concat_cp_element_group_300 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(300), clk => clk, reset => reset); --
    end block;
    -- CP-element group 301:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	197 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	330 
    -- CP-element group 301: marked-successors 
    -- CP-element group 301: 	195 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_final_index_sum_regn_sample_complete
      -- CP-element group 301: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_final_index_sum_regn_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_final_index_sum_regn_Sample/$exit
      -- 
    ack_1889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_845_index_offset_ack_0, ack => concat_CP_34_elements(301)); -- 
    -- CP-element group 302:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	300 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	298 
    -- CP-element group 302: marked-successors 
    -- CP-element group 302: 	300 
    -- CP-element group 302:  members (8) 
      -- CP-element group 302: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_base_plus_offset/sum_rename_req
      -- CP-element group 302: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_base_plus_offset/sum_rename_ack
      -- CP-element group 302: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_final_index_sum_regn_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_final_index_sum_regn_Update/ack
      -- CP-element group 302: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_base_plus_offset/$exit
      -- CP-element group 302: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_base_plus_offset/$entry
      -- CP-element group 302: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_offset_calculated
      -- CP-element group 302: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/array_obj_ref_845_root_address_calculated
      -- 
    ack_1894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_845_index_offset_ack_1, ack => concat_CP_34_elements(302)); -- 
    -- CP-element group 303:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	298 
    -- CP-element group 303: successors 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	298 
    -- CP-element group 303: 	300 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_846_request/$exit
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_846_request/ack
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_846_sample_completed_
      -- 
    ack_1904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_846_final_reg_ack_0, ack => concat_CP_34_elements(303)); -- 
    -- CP-element group 304:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	299 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304: marked-successors 
    -- CP-element group 304: 	299 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_846_complete/$exit
      -- CP-element group 304: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_846_complete/ack
      -- CP-element group 304: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/addr_of_846_update_completed_
      -- 
    ack_1909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_846_final_reg_ack_1, ack => concat_CP_34_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_850_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_850_Sample/req
      -- CP-element group 305: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_850_Sample/$entry
      -- 
    req_1917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(305), ack => W_ov_842_delayed_7_0_848_inst_req_0); -- 
    concat_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(304) & concat_CP_34_elements(307);
      gj_concat_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	308 
    -- CP-element group 306: 	319 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_850_Update/req
      -- CP-element group 306: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_850_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_850_update_start_
      -- 
    req_1922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(306), ack => W_ov_842_delayed_7_0_848_inst_req_1); -- 
    concat_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(308) & concat_CP_34_elements(319);
      gj_concat_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	299 
    -- CP-element group 307: 	305 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_850_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_850_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_850_Sample/$exit
      -- 
    ack_1918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ov_842_delayed_7_0_848_inst_ack_0, ack => concat_CP_34_elements(307)); -- 
    -- CP-element group 308:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	317 
    -- CP-element group 308: marked-successors 
    -- CP-element group 308: 	306 
    -- CP-element group 308:  members (19) 
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_word_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_base_address_resized
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_root_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_base_plus_offset/$entry
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_base_addr_resize/$entry
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_base_addr_resize/$exit
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_base_addr_resize/base_resize_req
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_base_addr_resize/base_resize_ack
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_base_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_850_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_850_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_850_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_word_addrgen/root_register_ack
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_word_addrgen/root_register_req
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_word_addrgen/$exit
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_word_addrgen/$entry
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_base_plus_offset/sum_rename_ack
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_base_plus_offset/sum_rename_req
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_base_plus_offset/$exit
      -- 
    ack_1923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ov_842_delayed_7_0_848_inst_ack_1, ack => concat_CP_34_elements(308)); -- 
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	254 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	311 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	311 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_853_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_853_Sample/req
      -- CP-element group 309: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_853_sample_start_
      -- 
    req_1931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(309), ack => W_cmp_844_delayed_12_0_851_inst_req_0); -- 
    concat_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(254) & concat_CP_34_elements(311);
      gj_concat_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	312 
    -- CP-element group 310: 	315 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_853_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_853_update_start_
      -- CP-element group 310: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_853_Update/req
      -- 
    req_1936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(310), ack => W_cmp_844_delayed_12_0_851_inst_req_1); -- 
    concat_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(312) & concat_CP_34_elements(315);
      gj_concat_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: successors 
    -- CP-element group 311: marked-successors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: 	250 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_853_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_853_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_853_Sample/ack
      -- 
    ack_1932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_cmp_844_delayed_12_0_851_inst_ack_0, ack => concat_CP_34_elements(311)); -- 
    -- CP-element group 312:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312: marked-successors 
    -- CP-element group 312: 	310 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_853_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_853_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/assign_stmt_853_Update/ack
      -- 
    ack_1937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_cmp_844_delayed_12_0_851_inst_ack_1, ack => concat_CP_34_elements(312)); -- 
    -- CP-element group 313:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: 	282 
    -- CP-element group 313: 	297 
    -- CP-element group 313: marked-predecessors 
    -- CP-element group 313: 	315 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	315 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/MUX_859_start/$entry
      -- CP-element group 313: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/MUX_859_sample_start_
      -- CP-element group 313: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/MUX_859_start/req
      -- 
    req_1945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(313), ack => MUX_859_inst_req_0); -- 
    concat_cp_element_group_313: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_313"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(312) & concat_CP_34_elements(282) & concat_CP_34_elements(297) & concat_CP_34_elements(315);
      gj_concat_cp_element_group_313 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(313), clk => clk, reset => reset); --
    end block;
    -- CP-element group 314:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: marked-predecessors 
    -- CP-element group 314: 	316 
    -- CP-element group 314: 	319 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	316 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/MUX_859_complete/$entry
      -- CP-element group 314: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/MUX_859_update_start_
      -- CP-element group 314: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/MUX_859_complete/req
      -- 
    req_1950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(314), ack => MUX_859_inst_req_1); -- 
    concat_cp_element_group_314: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_314"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(316) & concat_CP_34_elements(319);
      gj_concat_cp_element_group_314 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(314), clk => clk, reset => reset); --
    end block;
    -- CP-element group 315:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	313 
    -- CP-element group 315: successors 
    -- CP-element group 315: marked-successors 
    -- CP-element group 315: 	310 
    -- CP-element group 315: 	313 
    -- CP-element group 315: 	280 
    -- CP-element group 315: 	295 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/MUX_859_start/ack
      -- CP-element group 315: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/MUX_859_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/MUX_859_start/$exit
      -- 
    ack_1946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_859_inst_ack_0, ack => concat_CP_34_elements(315)); -- 
    -- CP-element group 316:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	314 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316: marked-successors 
    -- CP-element group 316: 	314 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/MUX_859_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/MUX_859_complete/$exit
      -- CP-element group 316: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/MUX_859_complete/ack
      -- 
    ack_1951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_859_inst_ack_1, ack => concat_CP_34_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	308 
    -- CP-element group 317: 	316 
    -- CP-element group 317: marked-predecessors 
    -- CP-element group 317: 	319 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	319 
    -- CP-element group 317:  members (9) 
      -- CP-element group 317: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Sample/word_access_start/word_0/rr
      -- CP-element group 317: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Sample/word_access_start/word_0/$entry
      -- CP-element group 317: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Sample/word_access_start/$entry
      -- CP-element group 317: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Sample/ptr_deref_855_Split/split_ack
      -- CP-element group 317: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Sample/ptr_deref_855_Split/split_req
      -- CP-element group 317: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Sample/ptr_deref_855_Split/$exit
      -- CP-element group 317: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Sample/ptr_deref_855_Split/$entry
      -- CP-element group 317: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Sample/$entry
      -- 
    rr_1989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(317), ack => ptr_deref_855_store_0_req_0); -- 
    concat_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(308) & concat_CP_34_elements(316) & concat_CP_34_elements(319);
      gj_concat_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: marked-predecessors 
    -- CP-element group 318: 	320 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	320 
    -- CP-element group 318:  members (5) 
      -- CP-element group 318: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_update_start_
      -- CP-element group 318: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Update/word_access_complete/word_0/cr
      -- CP-element group 318: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Update/word_access_complete/word_0/$entry
      -- CP-element group 318: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Update/word_access_complete/$entry
      -- CP-element group 318: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Update/$entry
      -- 
    cr_2000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(318), ack => ptr_deref_855_store_0_req_1); -- 
    concat_cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_318"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(320);
      gj_concat_cp_element_group_318 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 319:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	317 
    -- CP-element group 319: successors 
    -- CP-element group 319: marked-successors 
    -- CP-element group 319: 	314 
    -- CP-element group 319: 	317 
    -- CP-element group 319: 	306 
    -- CP-element group 319:  members (5) 
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Sample/word_access_start/word_0/ra
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Sample/word_access_start/word_0/$exit
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Sample/word_access_start/$exit
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Sample/$exit
      -- 
    ra_1990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_855_store_0_ack_0, ack => concat_CP_34_elements(319)); -- 
    -- CP-element group 320:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	318 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	330 
    -- CP-element group 320: marked-successors 
    -- CP-element group 320: 	318 
    -- CP-element group 320:  members (5) 
      -- CP-element group 320: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_update_completed_
      -- CP-element group 320: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Update/word_access_complete/word_0/ca
      -- CP-element group 320: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Update/word_access_complete/word_0/$exit
      -- CP-element group 320: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Update/word_access_complete/$exit
      -- CP-element group 320: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/ptr_deref_855_Update/$exit
      -- 
    ca_2001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_855_store_0_ack_1, ack => concat_CP_34_elements(320)); -- 
    -- CP-element group 321:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	188 
    -- CP-element group 321: marked-predecessors 
    -- CP-element group 321: 	323 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	323 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u16_u16_864_Sample/rr
      -- CP-element group 321: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u16_u16_864_Sample/$entry
      -- CP-element group 321: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u16_u16_864_sample_start_
      -- 
    rr_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(321), ack => SUB_u16_u16_864_inst_req_0); -- 
    concat_cp_element_group_321: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_321"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(323);
      gj_concat_cp_element_group_321 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(321), clk => clk, reset => reset); --
    end block;
    -- CP-element group 322:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	191 
    -- CP-element group 322: marked-predecessors 
    -- CP-element group 322: 	324 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u16_u16_864_Update/cr
      -- CP-element group 322: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u16_u16_864_Update/$entry
      -- CP-element group 322: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u16_u16_864_update_start_
      -- 
    cr_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(322), ack => SUB_u16_u16_864_inst_req_1); -- 
    concat_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(191) & concat_CP_34_elements(324);
      gj_concat_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	321 
    -- CP-element group 323: successors 
    -- CP-element group 323: marked-successors 
    -- CP-element group 323: 	321 
    -- CP-element group 323:  members (3) 
      -- CP-element group 323: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u16_u16_864_Sample/ra
      -- CP-element group 323: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u16_u16_864_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u16_u16_864_sample_completed_
      -- 
    ra_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_864_inst_ack_0, ack => concat_CP_34_elements(323)); -- 
    -- CP-element group 324:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	189 
    -- CP-element group 324: marked-successors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: 	249 
    -- CP-element group 324:  members (3) 
      -- CP-element group 324: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u16_u16_864_Update/ca
      -- CP-element group 324: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u16_u16_864_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u16_u16_864_update_completed_
      -- 
    ca_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_864_inst_ack_1, ack => concat_CP_34_elements(324)); -- 
    -- CP-element group 325:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	188 
    -- CP-element group 325: marked-predecessors 
    -- CP-element group 325: 	327 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	327 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u32_u32_903_sample_start_
      -- CP-element group 325: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u32_u32_903_Sample/rr
      -- CP-element group 325: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u32_u32_903_Sample/$entry
      -- 
    rr_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(325), ack => SUB_u32_u32_903_inst_req_0); -- 
    concat_cp_element_group_325: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_325"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(188) & concat_CP_34_elements(327);
      gj_concat_cp_element_group_325 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(325), clk => clk, reset => reset); --
    end block;
    -- CP-element group 326:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: marked-predecessors 
    -- CP-element group 326: 	328 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	328 
    -- CP-element group 326:  members (3) 
      -- CP-element group 326: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u32_u32_903_Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u32_u32_903_Update/cr
      -- CP-element group 326: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u32_u32_903_update_start_
      -- 
    cr_2028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(326), ack => SUB_u32_u32_903_inst_req_1); -- 
    concat_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(328);
      gj_concat_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: successors 
    -- CP-element group 327: marked-successors 
    -- CP-element group 327: 	325 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u32_u32_903_Sample/ra
      -- CP-element group 327: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u32_u32_903_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u32_u32_903_sample_completed_
      -- 
    ra_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_903_inst_ack_0, ack => concat_CP_34_elements(327)); -- 
    -- CP-element group 328:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	189 
    -- CP-element group 328: marked-successors 
    -- CP-element group 328: 	326 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u32_u32_903_Update/ca
      -- CP-element group 328: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u32_u32_903_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/SUB_u32_u32_903_update_completed_
      -- 
    ca_2029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_903_inst_ack_1, ack => concat_CP_34_elements(328)); -- 
    -- CP-element group 329:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	188 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	189 
    -- CP-element group 329:  members (1) 
      -- CP-element group 329: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group concat_CP_34_elements(329) is a control-delay.
    cp_element_329_delay: control_delay_element  generic map(name => " 329_delay", delay_value => 1)  port map(req => concat_CP_34_elements(188), ack => concat_CP_34_elements(329), clk => clk, reset =>reset);
    -- CP-element group 330:  join  transition  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	191 
    -- CP-element group 330: 	320 
    -- CP-element group 330: 	271 
    -- CP-element group 330: 	286 
    -- CP-element group 330: 	301 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	185 
    -- CP-element group 330:  members (1) 
      -- CP-element group 330: 	 branch_block_stmt_23/do_while_stmt_784/do_while_stmt_784_loop_body/$exit
      -- 
    concat_cp_element_group_330: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_330"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(191) & concat_CP_34_elements(320) & concat_CP_34_elements(271) & concat_CP_34_elements(286) & concat_CP_34_elements(301);
      gj_concat_cp_element_group_330 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(330), clk => clk, reset => reset); --
    end block;
    -- CP-element group 331:  transition  input  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	184 
    -- CP-element group 331: successors 
    -- CP-element group 331:  members (2) 
      -- CP-element group 331: 	 branch_block_stmt_23/do_while_stmt_784/loop_exit/$exit
      -- CP-element group 331: 	 branch_block_stmt_23/do_while_stmt_784/loop_exit/ack
      -- 
    ack_2034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_784_branch_ack_0, ack => concat_CP_34_elements(331)); -- 
    -- CP-element group 332:  transition  input  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	184 
    -- CP-element group 332: successors 
    -- CP-element group 332:  members (2) 
      -- CP-element group 332: 	 branch_block_stmt_23/do_while_stmt_784/loop_taken/$exit
      -- CP-element group 332: 	 branch_block_stmt_23/do_while_stmt_784/loop_taken/ack
      -- 
    ack_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_784_branch_ack_1, ack => concat_CP_34_elements(332)); -- 
    -- CP-element group 333:  transition  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	182 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	1 
    -- CP-element group 333:  members (1) 
      -- CP-element group 333: 	 branch_block_stmt_23/do_while_stmt_784/$exit
      -- 
    concat_CP_34_elements(333) <= concat_CP_34_elements(182);
    -- CP-element group 334:  transition  input  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	1 
    -- CP-element group 334: successors 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/call_stmt_917_Sample/$exit
      -- CP-element group 334: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/call_stmt_917_Sample/cra
      -- CP-element group 334: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/call_stmt_917_sample_completed_
      -- 
    cra_2051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_917_call_ack_0, ack => concat_CP_34_elements(334)); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	1 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	338 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/call_stmt_917_Update/$exit
      -- CP-element group 335: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/call_stmt_917_update_completed_
      -- CP-element group 335: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/call_stmt_917_Update/cca
      -- CP-element group 335: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_927_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_927_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_927_Sample/rr
      -- 
    cca_2056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_917_call_ack_1, ack => concat_CP_34_elements(335)); -- 
    rr_2078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(335), ack => type_cast_927_inst_req_0); -- 
    -- CP-element group 336:  transition  input  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	1 
    -- CP-element group 336: successors 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_922_Sample/$exit
      -- CP-element group 336: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_922_sample_completed_
      -- CP-element group 336: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_922_Sample/ra
      -- 
    ra_2065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_922_inst_ack_0, ack => concat_CP_34_elements(336)); -- 
    -- CP-element group 337:  fork  transition  input  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	1 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	340 
    -- CP-element group 337: 	343 
    -- CP-element group 337: 	346 
    -- CP-element group 337: 	349 
    -- CP-element group 337: 	352 
    -- CP-element group 337: 	355 
    -- CP-element group 337: 	358 
    -- CP-element group 337: 	361 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_922_update_completed_
      -- CP-element group 337: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_922_Update/$exit
      -- CP-element group 337: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_922_Update/ca
      -- 
    ca_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_922_inst_ack_1, ack => concat_CP_34_elements(337)); -- 
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	335 
    -- CP-element group 338: successors 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_927_sample_completed_
      -- CP-element group 338: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_927_Sample/$exit
      -- CP-element group 338: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_927_Sample/ra
      -- 
    ra_2079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_0, ack => concat_CP_34_elements(338)); -- 
    -- CP-element group 339:  fork  transition  input  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	1 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339: 	343 
    -- CP-element group 339: 	346 
    -- CP-element group 339: 	349 
    -- CP-element group 339: 	352 
    -- CP-element group 339: 	355 
    -- CP-element group 339: 	358 
    -- CP-element group 339: 	361 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_927_update_completed_
      -- CP-element group 339: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_927_Update/$exit
      -- CP-element group 339: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_927_Update/ca
      -- 
    ca_2084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_1, ack => concat_CP_34_elements(339)); -- 
    -- CP-element group 340:  join  transition  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	337 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_936_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_936_Sample/rr
      -- CP-element group 340: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_936_sample_start_
      -- 
    rr_2092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(340), ack => type_cast_936_inst_req_0); -- 
    concat_cp_element_group_340: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_340"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(337) & concat_CP_34_elements(339);
      gj_concat_cp_element_group_340 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(340), clk => clk, reset => reset); --
    end block;
    -- CP-element group 341:  transition  input  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_936_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_936_Sample/ra
      -- CP-element group 341: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_936_sample_completed_
      -- 
    ra_2093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_936_inst_ack_0, ack => concat_CP_34_elements(341)); -- 
    -- CP-element group 342:  transition  input  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	1 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	384 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_936_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_936_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_936_Update/ca
      -- 
    ca_2098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_936_inst_ack_1, ack => concat_CP_34_elements(342)); -- 
    -- CP-element group 343:  join  transition  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	337 
    -- CP-element group 343: 	339 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_946_sample_start_
      -- CP-element group 343: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_946_Sample/$entry
      -- CP-element group 343: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_946_Sample/rr
      -- 
    rr_2106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(343), ack => type_cast_946_inst_req_0); -- 
    concat_cp_element_group_343: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_343"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(337) & concat_CP_34_elements(339);
      gj_concat_cp_element_group_343 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(343), clk => clk, reset => reset); --
    end block;
    -- CP-element group 344:  transition  input  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_946_Sample/ra
      -- CP-element group 344: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_946_sample_completed_
      -- CP-element group 344: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_946_Sample/$exit
      -- 
    ra_2107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_946_inst_ack_0, ack => concat_CP_34_elements(344)); -- 
    -- CP-element group 345:  transition  input  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	1 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	381 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_946_update_completed_
      -- CP-element group 345: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_946_Update/ca
      -- CP-element group 345: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_946_Update/$exit
      -- 
    ca_2112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_946_inst_ack_1, ack => concat_CP_34_elements(345)); -- 
    -- CP-element group 346:  join  transition  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	337 
    -- CP-element group 346: 	339 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_956_Sample/rr
      -- CP-element group 346: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_956_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_956_sample_start_
      -- 
    rr_2120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(346), ack => type_cast_956_inst_req_0); -- 
    concat_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(337) & concat_CP_34_elements(339);
      gj_concat_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_956_Sample/ra
      -- CP-element group 347: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_956_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_956_sample_completed_
      -- 
    ra_2121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_956_inst_ack_0, ack => concat_CP_34_elements(347)); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	1 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	378 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_956_Update/ca
      -- CP-element group 348: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_956_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_956_update_completed_
      -- 
    ca_2126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_956_inst_ack_1, ack => concat_CP_34_elements(348)); -- 
    -- CP-element group 349:  join  transition  output  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	337 
    -- CP-element group 349: 	339 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	350 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_966_sample_start_
      -- CP-element group 349: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_966_Sample/$entry
      -- CP-element group 349: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_966_Sample/rr
      -- 
    rr_2134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(349), ack => type_cast_966_inst_req_0); -- 
    concat_cp_element_group_349: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_349"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(337) & concat_CP_34_elements(339);
      gj_concat_cp_element_group_349 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(349), clk => clk, reset => reset); --
    end block;
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	349 
    -- CP-element group 350: successors 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_966_sample_completed_
      -- CP-element group 350: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_966_Sample/$exit
      -- CP-element group 350: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_966_Sample/ra
      -- 
    ra_2135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_966_inst_ack_0, ack => concat_CP_34_elements(350)); -- 
    -- CP-element group 351:  transition  input  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	1 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	375 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_966_update_completed_
      -- CP-element group 351: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_966_Update/ca
      -- CP-element group 351: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_966_Update/$exit
      -- 
    ca_2140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_966_inst_ack_1, ack => concat_CP_34_elements(351)); -- 
    -- CP-element group 352:  join  transition  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	337 
    -- CP-element group 352: 	339 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_976_Sample/rr
      -- CP-element group 352: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_976_Sample/$entry
      -- CP-element group 352: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_976_sample_start_
      -- 
    rr_2148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(352), ack => type_cast_976_inst_req_0); -- 
    concat_cp_element_group_352: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_352"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(337) & concat_CP_34_elements(339);
      gj_concat_cp_element_group_352 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(352), clk => clk, reset => reset); --
    end block;
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_976_Sample/ra
      -- CP-element group 353: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_976_Sample/$exit
      -- CP-element group 353: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_976_sample_completed_
      -- 
    ra_2149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_976_inst_ack_0, ack => concat_CP_34_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	1 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	372 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_976_Update/ca
      -- CP-element group 354: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_976_Update/$exit
      -- CP-element group 354: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_976_update_completed_
      -- 
    ca_2154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_976_inst_ack_1, ack => concat_CP_34_elements(354)); -- 
    -- CP-element group 355:  join  transition  output  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	337 
    -- CP-element group 355: 	339 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_986_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_986_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_986_Sample/rr
      -- 
    rr_2162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(355), ack => type_cast_986_inst_req_0); -- 
    concat_cp_element_group_355: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_355"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(337) & concat_CP_34_elements(339);
      gj_concat_cp_element_group_355 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(355), clk => clk, reset => reset); --
    end block;
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_986_Sample/ra
      -- CP-element group 356: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_986_sample_completed_
      -- CP-element group 356: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_986_Sample/$exit
      -- 
    ra_2163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_986_inst_ack_0, ack => concat_CP_34_elements(356)); -- 
    -- CP-element group 357:  transition  input  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	1 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	369 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_986_update_completed_
      -- CP-element group 357: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_986_Update/ca
      -- CP-element group 357: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_986_Update/$exit
      -- 
    ca_2168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_986_inst_ack_1, ack => concat_CP_34_elements(357)); -- 
    -- CP-element group 358:  join  transition  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	337 
    -- CP-element group 358: 	339 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_996_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_996_Sample/rr
      -- CP-element group 358: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_996_Sample/$entry
      -- 
    rr_2176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(358), ack => type_cast_996_inst_req_0); -- 
    concat_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(337) & concat_CP_34_elements(339);
      gj_concat_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  transition  input  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_996_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_996_Sample/ra
      -- CP-element group 359: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_996_Sample/$exit
      -- 
    ra_2177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_996_inst_ack_0, ack => concat_CP_34_elements(359)); -- 
    -- CP-element group 360:  transition  input  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	1 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	366 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_996_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_996_Update/ca
      -- CP-element group 360: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_996_Update/$exit
      -- 
    ca_2182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_996_inst_ack_1, ack => concat_CP_34_elements(360)); -- 
    -- CP-element group 361:  join  transition  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	337 
    -- CP-element group 361: 	339 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_1006_Sample/rr
      -- CP-element group 361: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_1006_Sample/$entry
      -- CP-element group 361: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_1006_sample_start_
      -- 
    rr_2190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(361), ack => type_cast_1006_inst_req_0); -- 
    concat_cp_element_group_361: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_361"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(337) & concat_CP_34_elements(339);
      gj_concat_cp_element_group_361 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362:  members (3) 
      -- CP-element group 362: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_1006_Sample/ra
      -- CP-element group 362: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_1006_Sample/$exit
      -- CP-element group 362: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_1006_sample_completed_
      -- 
    ra_2191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1006_inst_ack_0, ack => concat_CP_34_elements(362)); -- 
    -- CP-element group 363:  transition  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	1 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1008_Sample/req
      -- CP-element group 363: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1008_Sample/$entry
      -- CP-element group 363: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1008_sample_start_
      -- CP-element group 363: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_1006_Update/ca
      -- CP-element group 363: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_1006_Update/$exit
      -- CP-element group 363: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/type_cast_1006_update_completed_
      -- 
    ca_2196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1006_inst_ack_1, ack => concat_CP_34_elements(363)); -- 
    req_2204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(363), ack => WPIPE_Concat_output_pipe_1008_inst_req_0); -- 
    -- CP-element group 364:  transition  input  output  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (6) 
      -- CP-element group 364: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1008_Update/req
      -- CP-element group 364: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1008_Update/$entry
      -- CP-element group 364: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1008_Sample/ack
      -- CP-element group 364: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1008_Sample/$exit
      -- CP-element group 364: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1008_update_start_
      -- CP-element group 364: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1008_sample_completed_
      -- 
    ack_2205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1008_inst_ack_0, ack => concat_CP_34_elements(364)); -- 
    req_2209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(364), ack => WPIPE_Concat_output_pipe_1008_inst_req_1); -- 
    -- CP-element group 365:  transition  input  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1008_Update/ack
      -- CP-element group 365: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1008_Update/$exit
      -- CP-element group 365: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1008_update_completed_
      -- 
    ack_2210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1008_inst_ack_1, ack => concat_CP_34_elements(365)); -- 
    -- CP-element group 366:  join  transition  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	360 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1011_Sample/req
      -- CP-element group 366: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1011_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1011_sample_start_
      -- 
    req_2218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(366), ack => WPIPE_Concat_output_pipe_1011_inst_req_0); -- 
    concat_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(360) & concat_CP_34_elements(365);
      gj_concat_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  transition  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (6) 
      -- CP-element group 367: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1011_Update/$entry
      -- CP-element group 367: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1011_Update/req
      -- CP-element group 367: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1011_Sample/ack
      -- CP-element group 367: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1011_Sample/$exit
      -- CP-element group 367: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1011_update_start_
      -- CP-element group 367: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1011_sample_completed_
      -- 
    ack_2219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1011_inst_ack_0, ack => concat_CP_34_elements(367)); -- 
    req_2223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(367), ack => WPIPE_Concat_output_pipe_1011_inst_req_1); -- 
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1011_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1011_Update/ack
      -- CP-element group 368: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1011_update_completed_
      -- 
    ack_2224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1011_inst_ack_1, ack => concat_CP_34_elements(368)); -- 
    -- CP-element group 369:  join  transition  output  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	357 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1014_Sample/req
      -- CP-element group 369: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1014_Sample/$entry
      -- CP-element group 369: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1014_sample_start_
      -- 
    req_2232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(369), ack => WPIPE_Concat_output_pipe_1014_inst_req_0); -- 
    concat_cp_element_group_369: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_369"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(357) & concat_CP_34_elements(368);
      gj_concat_cp_element_group_369 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(369), clk => clk, reset => reset); --
    end block;
    -- CP-element group 370:  transition  input  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (6) 
      -- CP-element group 370: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1014_Update/req
      -- CP-element group 370: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1014_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1014_Sample/ack
      -- CP-element group 370: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1014_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1014_update_start_
      -- CP-element group 370: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1014_sample_completed_
      -- 
    ack_2233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1014_inst_ack_0, ack => concat_CP_34_elements(370)); -- 
    req_2237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(370), ack => WPIPE_Concat_output_pipe_1014_inst_req_1); -- 
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1014_Update/ack
      -- CP-element group 371: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1014_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1014_update_completed_
      -- 
    ack_2238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1014_inst_ack_1, ack => concat_CP_34_elements(371)); -- 
    -- CP-element group 372:  join  transition  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	354 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1017_Sample/req
      -- CP-element group 372: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1017_Sample/$entry
      -- CP-element group 372: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1017_sample_start_
      -- 
    req_2246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(372), ack => WPIPE_Concat_output_pipe_1017_inst_req_0); -- 
    concat_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(354) & concat_CP_34_elements(371);
      gj_concat_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  transition  input  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (6) 
      -- CP-element group 373: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1017_Update/req
      -- CP-element group 373: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1017_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1017_Sample/ack
      -- CP-element group 373: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1017_Sample/$exit
      -- CP-element group 373: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1017_update_start_
      -- CP-element group 373: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1017_sample_completed_
      -- 
    ack_2247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1017_inst_ack_0, ack => concat_CP_34_elements(373)); -- 
    req_2251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(373), ack => WPIPE_Concat_output_pipe_1017_inst_req_1); -- 
    -- CP-element group 374:  transition  input  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1017_Update/ack
      -- CP-element group 374: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1017_Update/$exit
      -- CP-element group 374: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1017_update_completed_
      -- 
    ack_2252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1017_inst_ack_1, ack => concat_CP_34_elements(374)); -- 
    -- CP-element group 375:  join  transition  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	351 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1020_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1020_Sample/req
      -- CP-element group 375: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1020_Sample/$entry
      -- 
    req_2260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(375), ack => WPIPE_Concat_output_pipe_1020_inst_req_0); -- 
    concat_cp_element_group_375: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_375"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(351) & concat_CP_34_elements(374);
      gj_concat_cp_element_group_375 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(375), clk => clk, reset => reset); --
    end block;
    -- CP-element group 376:  transition  input  output  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (6) 
      -- CP-element group 376: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1020_Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1020_Update/req
      -- CP-element group 376: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1020_Sample/ack
      -- CP-element group 376: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1020_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1020_update_start_
      -- CP-element group 376: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1020_sample_completed_
      -- 
    ack_2261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1020_inst_ack_0, ack => concat_CP_34_elements(376)); -- 
    req_2265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(376), ack => WPIPE_Concat_output_pipe_1020_inst_req_1); -- 
    -- CP-element group 377:  transition  input  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1020_Update/$exit
      -- CP-element group 377: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1020_Update/ack
      -- CP-element group 377: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1020_update_completed_
      -- 
    ack_2266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1020_inst_ack_1, ack => concat_CP_34_elements(377)); -- 
    -- CP-element group 378:  join  transition  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	348 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1023_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1023_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1023_Sample/req
      -- 
    req_2274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(378), ack => WPIPE_Concat_output_pipe_1023_inst_req_0); -- 
    concat_cp_element_group_378: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_378"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(348) & concat_CP_34_elements(377);
      gj_concat_cp_element_group_378 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(378), clk => clk, reset => reset); --
    end block;
    -- CP-element group 379:  transition  input  output  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379:  members (6) 
      -- CP-element group 379: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1023_Update/req
      -- CP-element group 379: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1023_sample_completed_
      -- CP-element group 379: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1023_Sample/$exit
      -- CP-element group 379: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1023_Update/$entry
      -- CP-element group 379: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1023_update_start_
      -- CP-element group 379: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1023_Sample/ack
      -- 
    ack_2275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1023_inst_ack_0, ack => concat_CP_34_elements(379)); -- 
    req_2279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(379), ack => WPIPE_Concat_output_pipe_1023_inst_req_1); -- 
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	379 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	381 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1023_update_completed_
      -- CP-element group 380: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1023_Update/$exit
      -- CP-element group 380: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1023_Update/ack
      -- 
    ack_2280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1023_inst_ack_1, ack => concat_CP_34_elements(380)); -- 
    -- CP-element group 381:  join  transition  output  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	345 
    -- CP-element group 381: 	380 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1026_sample_start_
      -- CP-element group 381: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1026_Sample/$entry
      -- CP-element group 381: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1026_Sample/req
      -- 
    req_2288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(381), ack => WPIPE_Concat_output_pipe_1026_inst_req_0); -- 
    concat_cp_element_group_381: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_381"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(345) & concat_CP_34_elements(380);
      gj_concat_cp_element_group_381 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(381), clk => clk, reset => reset); --
    end block;
    -- CP-element group 382:  transition  input  output  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382:  members (6) 
      -- CP-element group 382: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1026_sample_completed_
      -- CP-element group 382: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1026_update_start_
      -- CP-element group 382: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1026_Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1026_Sample/ack
      -- CP-element group 382: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1026_Update/$entry
      -- CP-element group 382: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1026_Update/req
      -- 
    ack_2289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1026_inst_ack_0, ack => concat_CP_34_elements(382)); -- 
    req_2293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(382), ack => WPIPE_Concat_output_pipe_1026_inst_req_1); -- 
    -- CP-element group 383:  transition  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	382 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1026_update_completed_
      -- CP-element group 383: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1026_Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1026_Update/ack
      -- 
    ack_2294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1026_inst_ack_1, ack => concat_CP_34_elements(383)); -- 
    -- CP-element group 384:  join  transition  output  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	342 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1029_sample_start_
      -- CP-element group 384: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1029_Sample/$entry
      -- CP-element group 384: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1029_Sample/req
      -- 
    req_2302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(384), ack => WPIPE_Concat_output_pipe_1029_inst_req_0); -- 
    concat_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(342) & concat_CP_34_elements(383);
      gj_concat_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  transition  input  output  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (6) 
      -- CP-element group 385: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1029_sample_completed_
      -- CP-element group 385: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1029_update_start_
      -- CP-element group 385: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1029_Sample/$exit
      -- CP-element group 385: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1029_Sample/ack
      -- CP-element group 385: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1029_Update/$entry
      -- CP-element group 385: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1029_Update/req
      -- 
    ack_2303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1029_inst_ack_0, ack => concat_CP_34_elements(385)); -- 
    req_2307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(385), ack => WPIPE_Concat_output_pipe_1029_inst_req_1); -- 
    -- CP-element group 386:  branch  transition  place  input  output  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	387 
    -- CP-element group 386: 	388 
    -- CP-element group 386:  members (17) 
      -- CP-element group 386: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031__exit__
      -- CP-element group 386: 	 branch_block_stmt_23/assign_stmt_1038__entry__
      -- CP-element group 386: 	 branch_block_stmt_23/assign_stmt_1038__exit__
      -- CP-element group 386: 	 branch_block_stmt_23/if_stmt_1039__entry__
      -- CP-element group 386: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/$exit
      -- CP-element group 386: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1029_update_completed_
      -- CP-element group 386: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1029_Update/$exit
      -- CP-element group 386: 	 branch_block_stmt_23/call_stmt_917_to_assign_stmt_1031/WPIPE_Concat_output_pipe_1029_Update/ack
      -- CP-element group 386: 	 branch_block_stmt_23/assign_stmt_1038/$entry
      -- CP-element group 386: 	 branch_block_stmt_23/assign_stmt_1038/$exit
      -- CP-element group 386: 	 branch_block_stmt_23/if_stmt_1039_dead_link/$entry
      -- CP-element group 386: 	 branch_block_stmt_23/if_stmt_1039_eval_test/$entry
      -- CP-element group 386: 	 branch_block_stmt_23/if_stmt_1039_eval_test/$exit
      -- CP-element group 386: 	 branch_block_stmt_23/if_stmt_1039_eval_test/branch_req
      -- CP-element group 386: 	 branch_block_stmt_23/R_cmp381460_1040_place
      -- CP-element group 386: 	 branch_block_stmt_23/if_stmt_1039_if_link/$entry
      -- CP-element group 386: 	 branch_block_stmt_23/if_stmt_1039_else_link/$entry
      -- 
    ack_2308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1029_inst_ack_1, ack => concat_CP_34_elements(386)); -- 
    branch_req_2319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(386), ack => if_stmt_1039_branch_req_0); -- 
    -- CP-element group 387:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	386 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	389 
    -- CP-element group 387: 	390 
    -- CP-element group 387:  members (18) 
      -- CP-element group 387: 	 branch_block_stmt_23/merge_stmt_1045__exit__
      -- CP-element group 387: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074__entry__
      -- CP-element group 387: 	 branch_block_stmt_23/merge_stmt_1045_PhiReqMerge
      -- CP-element group 387: 	 branch_block_stmt_23/if_stmt_1039_if_link/$exit
      -- CP-element group 387: 	 branch_block_stmt_23/if_stmt_1039_if_link/if_choice_transition
      -- CP-element group 387: 	 branch_block_stmt_23/whilex_xend_bbx_xnph
      -- CP-element group 387: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/$entry
      -- CP-element group 387: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/type_cast_1060_sample_start_
      -- CP-element group 387: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/type_cast_1060_update_start_
      -- CP-element group 387: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/type_cast_1060_Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/type_cast_1060_Sample/rr
      -- CP-element group 387: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/type_cast_1060_Update/$entry
      -- CP-element group 387: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/type_cast_1060_Update/cr
      -- CP-element group 387: 	 branch_block_stmt_23/merge_stmt_1045_PhiAck/dummy
      -- CP-element group 387: 	 branch_block_stmt_23/merge_stmt_1045_PhiAck/$exit
      -- CP-element group 387: 	 branch_block_stmt_23/merge_stmt_1045_PhiAck/$entry
      -- CP-element group 387: 	 branch_block_stmt_23/whilex_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 387: 	 branch_block_stmt_23/whilex_xend_bbx_xnph_PhiReq/$entry
      -- 
    if_choice_transition_2324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1039_branch_ack_1, ack => concat_CP_34_elements(387)); -- 
    rr_2341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(387), ack => type_cast_1060_inst_req_0); -- 
    cr_2346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(387), ack => type_cast_1060_inst_req_1); -- 
    -- CP-element group 388:  transition  place  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	386 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	459 
    -- CP-element group 388:  members (5) 
      -- CP-element group 388: 	 branch_block_stmt_23/if_stmt_1039_else_link/$exit
      -- CP-element group 388: 	 branch_block_stmt_23/if_stmt_1039_else_link/else_choice_transition
      -- CP-element group 388: 	 branch_block_stmt_23/whilex_xend_forx_xend456
      -- CP-element group 388: 	 branch_block_stmt_23/whilex_xend_forx_xend456_PhiReq/$exit
      -- CP-element group 388: 	 branch_block_stmt_23/whilex_xend_forx_xend456_PhiReq/$entry
      -- 
    else_choice_transition_2328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1039_branch_ack_0, ack => concat_CP_34_elements(388)); -- 
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	387 
    -- CP-element group 389: successors 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/type_cast_1060_sample_completed_
      -- CP-element group 389: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/type_cast_1060_Sample/$exit
      -- CP-element group 389: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/type_cast_1060_Sample/ra
      -- 
    ra_2342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1060_inst_ack_0, ack => concat_CP_34_elements(389)); -- 
    -- CP-element group 390:  transition  place  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	387 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	453 
    -- CP-element group 390:  members (9) 
      -- CP-element group 390: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074__exit__
      -- CP-element group 390: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383
      -- CP-element group 390: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/$exit
      -- CP-element group 390: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/type_cast_1060_update_completed_
      -- CP-element group 390: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/type_cast_1060_Update/$exit
      -- CP-element group 390: 	 branch_block_stmt_23/assign_stmt_1051_to_assign_stmt_1074/type_cast_1060_Update/ca
      -- CP-element group 390: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/$entry
      -- CP-element group 390: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/phi_stmt_1077/$entry
      -- CP-element group 390: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/$entry
      -- 
    ca_2347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1060_inst_ack_1, ack => concat_CP_34_elements(390)); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	458 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	436 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_final_index_sum_regn_sample_complete
      -- CP-element group 391: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_final_index_sum_regn_Sample/$exit
      -- CP-element group 391: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_final_index_sum_regn_Sample/ack
      -- 
    ack_2376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1089_index_offset_ack_0, ack => concat_CP_34_elements(391)); -- 
    -- CP-element group 392:  transition  input  output  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	458 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	393 
    -- CP-element group 392:  members (11) 
      -- CP-element group 392: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/addr_of_1090_sample_start_
      -- CP-element group 392: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_root_address_calculated
      -- CP-element group 392: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_offset_calculated
      -- CP-element group 392: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_final_index_sum_regn_Update/$exit
      -- CP-element group 392: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_final_index_sum_regn_Update/ack
      -- CP-element group 392: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_base_plus_offset/$entry
      -- CP-element group 392: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_base_plus_offset/$exit
      -- CP-element group 392: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_base_plus_offset/sum_rename_req
      -- CP-element group 392: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_base_plus_offset/sum_rename_ack
      -- CP-element group 392: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/addr_of_1090_request/$entry
      -- CP-element group 392: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/addr_of_1090_request/req
      -- 
    ack_2381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1089_index_offset_ack_1, ack => concat_CP_34_elements(392)); -- 
    req_2390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(392), ack => addr_of_1090_final_reg_req_0); -- 
    -- CP-element group 393:  transition  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	392 
    -- CP-element group 393: successors 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/addr_of_1090_sample_completed_
      -- CP-element group 393: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/addr_of_1090_request/$exit
      -- CP-element group 393: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/addr_of_1090_request/ack
      -- 
    ack_2391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1090_final_reg_ack_0, ack => concat_CP_34_elements(393)); -- 
    -- CP-element group 394:  join  fork  transition  input  output  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	458 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (24) 
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/addr_of_1090_update_completed_
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/addr_of_1090_complete/$exit
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/addr_of_1090_complete/ack
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_sample_start_
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_base_address_calculated
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_word_address_calculated
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_root_address_calculated
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_base_address_resized
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_base_addr_resize/$entry
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_base_addr_resize/$exit
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_base_addr_resize/base_resize_req
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_base_addr_resize/base_resize_ack
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_base_plus_offset/$entry
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_base_plus_offset/$exit
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_base_plus_offset/sum_rename_req
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_base_plus_offset/sum_rename_ack
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_word_addrgen/$entry
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_word_addrgen/$exit
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_word_addrgen/root_register_req
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_word_addrgen/root_register_ack
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Sample/$entry
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Sample/word_access_start/$entry
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Sample/word_access_start/word_0/$entry
      -- CP-element group 394: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Sample/word_access_start/word_0/rr
      -- 
    ack_2396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1090_final_reg_ack_1, ack => concat_CP_34_elements(394)); -- 
    rr_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(394), ack => ptr_deref_1094_load_0_req_0); -- 
    -- CP-element group 395:  transition  input  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395:  members (5) 
      -- CP-element group 395: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_sample_completed_
      -- CP-element group 395: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Sample/$exit
      -- CP-element group 395: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Sample/word_access_start/$exit
      -- CP-element group 395: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Sample/word_access_start/word_0/$exit
      -- CP-element group 395: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Sample/word_access_start/word_0/ra
      -- 
    ra_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1094_load_0_ack_0, ack => concat_CP_34_elements(395)); -- 
    -- CP-element group 396:  fork  transition  input  output  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	458 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396: 	399 
    -- CP-element group 396: 	401 
    -- CP-element group 396: 	403 
    -- CP-element group 396: 	405 
    -- CP-element group 396: 	407 
    -- CP-element group 396: 	409 
    -- CP-element group 396: 	411 
    -- CP-element group 396:  members (33) 
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_update_completed_
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Update/$exit
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Update/word_access_complete/$exit
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Update/word_access_complete/word_0/$exit
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Update/word_access_complete/word_0/ca
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Update/ptr_deref_1094_Merge/$entry
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Update/ptr_deref_1094_Merge/$exit
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Update/ptr_deref_1094_Merge/merge_req
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Update/ptr_deref_1094_Merge/merge_ack
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1098_sample_start_
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1098_Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1098_Sample/rr
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1108_sample_start_
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1108_Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1108_Sample/rr
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1118_sample_start_
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1118_Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1118_Sample/rr
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1128_sample_start_
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1128_Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1128_Sample/rr
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1138_sample_start_
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1138_Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1138_Sample/rr
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1148_sample_start_
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1148_Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1148_Sample/rr
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1158_sample_start_
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1158_Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1158_Sample/rr
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1168_sample_start_
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1168_Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1168_Sample/rr
      -- 
    ca_2441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1094_load_0_ack_1, ack => concat_CP_34_elements(396)); -- 
    rr_2454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(396), ack => type_cast_1098_inst_req_0); -- 
    rr_2468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(396), ack => type_cast_1108_inst_req_0); -- 
    rr_2482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(396), ack => type_cast_1118_inst_req_0); -- 
    rr_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(396), ack => type_cast_1128_inst_req_0); -- 
    rr_2510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(396), ack => type_cast_1138_inst_req_0); -- 
    rr_2524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(396), ack => type_cast_1148_inst_req_0); -- 
    rr_2538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(396), ack => type_cast_1158_inst_req_0); -- 
    rr_2552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(396), ack => type_cast_1168_inst_req_0); -- 
    -- CP-element group 397:  transition  input  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1098_sample_completed_
      -- CP-element group 397: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1098_Sample/$exit
      -- CP-element group 397: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1098_Sample/ra
      -- 
    ra_2455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1098_inst_ack_0, ack => concat_CP_34_elements(397)); -- 
    -- CP-element group 398:  transition  input  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	458 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	433 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1098_update_completed_
      -- CP-element group 398: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1098_Update/$exit
      -- CP-element group 398: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1098_Update/ca
      -- 
    ca_2460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1098_inst_ack_1, ack => concat_CP_34_elements(398)); -- 
    -- CP-element group 399:  transition  input  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	396 
    -- CP-element group 399: successors 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1108_sample_completed_
      -- CP-element group 399: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1108_Sample/$exit
      -- CP-element group 399: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1108_Sample/ra
      -- 
    ra_2469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1108_inst_ack_0, ack => concat_CP_34_elements(399)); -- 
    -- CP-element group 400:  transition  input  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	458 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	430 
    -- CP-element group 400:  members (3) 
      -- CP-element group 400: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1108_update_completed_
      -- CP-element group 400: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1108_Update/$exit
      -- CP-element group 400: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1108_Update/ca
      -- 
    ca_2474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1108_inst_ack_1, ack => concat_CP_34_elements(400)); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	396 
    -- CP-element group 401: successors 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1118_sample_completed_
      -- CP-element group 401: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1118_Sample/$exit
      -- CP-element group 401: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1118_Sample/ra
      -- 
    ra_2483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1118_inst_ack_0, ack => concat_CP_34_elements(401)); -- 
    -- CP-element group 402:  transition  input  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	458 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	427 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1118_update_completed_
      -- CP-element group 402: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1118_Update/$exit
      -- CP-element group 402: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1118_Update/ca
      -- 
    ca_2488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1118_inst_ack_1, ack => concat_CP_34_elements(402)); -- 
    -- CP-element group 403:  transition  input  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	396 
    -- CP-element group 403: successors 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1128_sample_completed_
      -- CP-element group 403: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1128_Sample/$exit
      -- CP-element group 403: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1128_Sample/ra
      -- 
    ra_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1128_inst_ack_0, ack => concat_CP_34_elements(403)); -- 
    -- CP-element group 404:  transition  input  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	458 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	424 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1128_update_completed_
      -- CP-element group 404: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1128_Update/$exit
      -- CP-element group 404: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1128_Update/ca
      -- 
    ca_2502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1128_inst_ack_1, ack => concat_CP_34_elements(404)); -- 
    -- CP-element group 405:  transition  input  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	396 
    -- CP-element group 405: successors 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1138_sample_completed_
      -- CP-element group 405: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1138_Sample/$exit
      -- CP-element group 405: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1138_Sample/ra
      -- 
    ra_2511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1138_inst_ack_0, ack => concat_CP_34_elements(405)); -- 
    -- CP-element group 406:  transition  input  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	458 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	421 
    -- CP-element group 406:  members (3) 
      -- CP-element group 406: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1138_update_completed_
      -- CP-element group 406: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1138_Update/$exit
      -- CP-element group 406: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1138_Update/ca
      -- 
    ca_2516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1138_inst_ack_1, ack => concat_CP_34_elements(406)); -- 
    -- CP-element group 407:  transition  input  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	396 
    -- CP-element group 407: successors 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1148_sample_completed_
      -- CP-element group 407: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1148_Sample/$exit
      -- CP-element group 407: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1148_Sample/ra
      -- 
    ra_2525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1148_inst_ack_0, ack => concat_CP_34_elements(407)); -- 
    -- CP-element group 408:  transition  input  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	458 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	418 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1148_update_completed_
      -- CP-element group 408: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1148_Update/$exit
      -- CP-element group 408: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1148_Update/ca
      -- 
    ca_2530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1148_inst_ack_1, ack => concat_CP_34_elements(408)); -- 
    -- CP-element group 409:  transition  input  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	396 
    -- CP-element group 409: successors 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1158_sample_completed_
      -- CP-element group 409: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1158_Sample/$exit
      -- CP-element group 409: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1158_Sample/ra
      -- 
    ra_2539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1158_inst_ack_0, ack => concat_CP_34_elements(409)); -- 
    -- CP-element group 410:  transition  input  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	458 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	415 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1158_update_completed_
      -- CP-element group 410: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1158_Update/$exit
      -- CP-element group 410: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1158_Update/ca
      -- 
    ca_2544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1158_inst_ack_1, ack => concat_CP_34_elements(410)); -- 
    -- CP-element group 411:  transition  input  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	396 
    -- CP-element group 411: successors 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1168_sample_completed_
      -- CP-element group 411: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1168_Sample/$exit
      -- CP-element group 411: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1168_Sample/ra
      -- 
    ra_2553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1168_inst_ack_0, ack => concat_CP_34_elements(411)); -- 
    -- CP-element group 412:  transition  input  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	458 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (6) 
      -- CP-element group 412: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1168_update_completed_
      -- CP-element group 412: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1168_Update/$exit
      -- CP-element group 412: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1168_Update/ca
      -- CP-element group 412: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1170_sample_start_
      -- CP-element group 412: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1170_Sample/$entry
      -- CP-element group 412: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1170_Sample/req
      -- 
    ca_2558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1168_inst_ack_1, ack => concat_CP_34_elements(412)); -- 
    req_2566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(412), ack => WPIPE_Concat_output_pipe_1170_inst_req_0); -- 
    -- CP-element group 413:  transition  input  output  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (6) 
      -- CP-element group 413: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1170_sample_completed_
      -- CP-element group 413: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1170_update_start_
      -- CP-element group 413: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1170_Sample/$exit
      -- CP-element group 413: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1170_Sample/ack
      -- CP-element group 413: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1170_Update/$entry
      -- CP-element group 413: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1170_Update/req
      -- 
    ack_2567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1170_inst_ack_0, ack => concat_CP_34_elements(413)); -- 
    req_2571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(413), ack => WPIPE_Concat_output_pipe_1170_inst_req_1); -- 
    -- CP-element group 414:  transition  input  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1170_update_completed_
      -- CP-element group 414: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1170_Update/$exit
      -- CP-element group 414: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1170_Update/ack
      -- 
    ack_2572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1170_inst_ack_1, ack => concat_CP_34_elements(414)); -- 
    -- CP-element group 415:  join  transition  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	410 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1173_sample_start_
      -- CP-element group 415: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1173_Sample/$entry
      -- CP-element group 415: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1173_Sample/req
      -- 
    req_2580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(415), ack => WPIPE_Concat_output_pipe_1173_inst_req_0); -- 
    concat_cp_element_group_415: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_415"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(410) & concat_CP_34_elements(414);
      gj_concat_cp_element_group_415 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(415), clk => clk, reset => reset); --
    end block;
    -- CP-element group 416:  transition  input  output  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416:  members (6) 
      -- CP-element group 416: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1173_sample_completed_
      -- CP-element group 416: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1173_update_start_
      -- CP-element group 416: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1173_Sample/$exit
      -- CP-element group 416: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1173_Sample/ack
      -- CP-element group 416: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1173_Update/$entry
      -- CP-element group 416: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1173_Update/req
      -- 
    ack_2581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1173_inst_ack_0, ack => concat_CP_34_elements(416)); -- 
    req_2585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(416), ack => WPIPE_Concat_output_pipe_1173_inst_req_1); -- 
    -- CP-element group 417:  transition  input  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	418 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1173_update_completed_
      -- CP-element group 417: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1173_Update/$exit
      -- CP-element group 417: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1173_Update/ack
      -- 
    ack_2586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1173_inst_ack_1, ack => concat_CP_34_elements(417)); -- 
    -- CP-element group 418:  join  transition  output  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	408 
    -- CP-element group 418: 	417 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	419 
    -- CP-element group 418:  members (3) 
      -- CP-element group 418: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1176_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1176_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1176_Sample/req
      -- 
    req_2594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(418), ack => WPIPE_Concat_output_pipe_1176_inst_req_0); -- 
    concat_cp_element_group_418: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_418"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(408) & concat_CP_34_elements(417);
      gj_concat_cp_element_group_418 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(418), clk => clk, reset => reset); --
    end block;
    -- CP-element group 419:  transition  input  output  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	418 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	420 
    -- CP-element group 419:  members (6) 
      -- CP-element group 419: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1176_sample_completed_
      -- CP-element group 419: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1176_update_start_
      -- CP-element group 419: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1176_Sample/$exit
      -- CP-element group 419: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1176_Sample/ack
      -- CP-element group 419: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1176_Update/$entry
      -- CP-element group 419: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1176_Update/req
      -- 
    ack_2595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1176_inst_ack_0, ack => concat_CP_34_elements(419)); -- 
    req_2599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(419), ack => WPIPE_Concat_output_pipe_1176_inst_req_1); -- 
    -- CP-element group 420:  transition  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	419 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	421 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1176_update_completed_
      -- CP-element group 420: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1176_Update/$exit
      -- CP-element group 420: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1176_Update/ack
      -- 
    ack_2600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1176_inst_ack_1, ack => concat_CP_34_elements(420)); -- 
    -- CP-element group 421:  join  transition  output  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	406 
    -- CP-element group 421: 	420 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	422 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1179_sample_start_
      -- CP-element group 421: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1179_Sample/$entry
      -- CP-element group 421: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1179_Sample/req
      -- 
    req_2608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(421), ack => WPIPE_Concat_output_pipe_1179_inst_req_0); -- 
    concat_cp_element_group_421: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_421"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(406) & concat_CP_34_elements(420);
      gj_concat_cp_element_group_421 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(421), clk => clk, reset => reset); --
    end block;
    -- CP-element group 422:  transition  input  output  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	421 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (6) 
      -- CP-element group 422: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1179_sample_completed_
      -- CP-element group 422: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1179_update_start_
      -- CP-element group 422: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1179_Sample/$exit
      -- CP-element group 422: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1179_Sample/ack
      -- CP-element group 422: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1179_Update/$entry
      -- CP-element group 422: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1179_Update/req
      -- 
    ack_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1179_inst_ack_0, ack => concat_CP_34_elements(422)); -- 
    req_2613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(422), ack => WPIPE_Concat_output_pipe_1179_inst_req_1); -- 
    -- CP-element group 423:  transition  input  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1179_update_completed_
      -- CP-element group 423: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1179_Update/$exit
      -- CP-element group 423: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1179_Update/ack
      -- 
    ack_2614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1179_inst_ack_1, ack => concat_CP_34_elements(423)); -- 
    -- CP-element group 424:  join  transition  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	404 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	425 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1182_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1182_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1182_Sample/req
      -- 
    req_2622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(424), ack => WPIPE_Concat_output_pipe_1182_inst_req_0); -- 
    concat_cp_element_group_424: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_424"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(404) & concat_CP_34_elements(423);
      gj_concat_cp_element_group_424 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(424), clk => clk, reset => reset); --
    end block;
    -- CP-element group 425:  transition  input  output  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	424 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425:  members (6) 
      -- CP-element group 425: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1182_sample_completed_
      -- CP-element group 425: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1182_update_start_
      -- CP-element group 425: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1182_Sample/$exit
      -- CP-element group 425: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1182_Sample/ack
      -- CP-element group 425: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1182_Update/$entry
      -- CP-element group 425: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1182_Update/req
      -- 
    ack_2623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1182_inst_ack_0, ack => concat_CP_34_elements(425)); -- 
    req_2627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(425), ack => WPIPE_Concat_output_pipe_1182_inst_req_1); -- 
    -- CP-element group 426:  transition  input  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426:  members (3) 
      -- CP-element group 426: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1182_update_completed_
      -- CP-element group 426: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1182_Update/$exit
      -- CP-element group 426: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1182_Update/ack
      -- 
    ack_2628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1182_inst_ack_1, ack => concat_CP_34_elements(426)); -- 
    -- CP-element group 427:  join  transition  output  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	402 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1185_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1185_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1185_Sample/req
      -- 
    req_2636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(427), ack => WPIPE_Concat_output_pipe_1185_inst_req_0); -- 
    concat_cp_element_group_427: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_427"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(402) & concat_CP_34_elements(426);
      gj_concat_cp_element_group_427 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(427), clk => clk, reset => reset); --
    end block;
    -- CP-element group 428:  transition  input  output  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	429 
    -- CP-element group 428:  members (6) 
      -- CP-element group 428: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1185_sample_completed_
      -- CP-element group 428: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1185_update_start_
      -- CP-element group 428: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1185_Sample/$exit
      -- CP-element group 428: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1185_Sample/ack
      -- CP-element group 428: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1185_Update/$entry
      -- CP-element group 428: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1185_Update/req
      -- 
    ack_2637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1185_inst_ack_0, ack => concat_CP_34_elements(428)); -- 
    req_2641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(428), ack => WPIPE_Concat_output_pipe_1185_inst_req_1); -- 
    -- CP-element group 429:  transition  input  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	428 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	430 
    -- CP-element group 429:  members (3) 
      -- CP-element group 429: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1185_update_completed_
      -- CP-element group 429: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1185_Update/$exit
      -- CP-element group 429: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1185_Update/ack
      -- 
    ack_2642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1185_inst_ack_1, ack => concat_CP_34_elements(429)); -- 
    -- CP-element group 430:  join  transition  output  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	400 
    -- CP-element group 430: 	429 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	431 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1188_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1188_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1188_Sample/req
      -- 
    req_2650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(430), ack => WPIPE_Concat_output_pipe_1188_inst_req_0); -- 
    concat_cp_element_group_430: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_430"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(400) & concat_CP_34_elements(429);
      gj_concat_cp_element_group_430 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(430), clk => clk, reset => reset); --
    end block;
    -- CP-element group 431:  transition  input  output  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	430 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	432 
    -- CP-element group 431:  members (6) 
      -- CP-element group 431: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1188_sample_completed_
      -- CP-element group 431: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1188_update_start_
      -- CP-element group 431: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1188_Sample/$exit
      -- CP-element group 431: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1188_Sample/ack
      -- CP-element group 431: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1188_Update/$entry
      -- CP-element group 431: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1188_Update/req
      -- 
    ack_2651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1188_inst_ack_0, ack => concat_CP_34_elements(431)); -- 
    req_2655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(431), ack => WPIPE_Concat_output_pipe_1188_inst_req_1); -- 
    -- CP-element group 432:  transition  input  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	431 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	433 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1188_update_completed_
      -- CP-element group 432: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1188_Update/$exit
      -- CP-element group 432: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1188_Update/ack
      -- 
    ack_2656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1188_inst_ack_1, ack => concat_CP_34_elements(432)); -- 
    -- CP-element group 433:  join  transition  output  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	398 
    -- CP-element group 433: 	432 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	434 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1191_sample_start_
      -- CP-element group 433: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1191_Sample/$entry
      -- CP-element group 433: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1191_Sample/req
      -- 
    req_2664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(433), ack => WPIPE_Concat_output_pipe_1191_inst_req_0); -- 
    concat_cp_element_group_433: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_433"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(398) & concat_CP_34_elements(432);
      gj_concat_cp_element_group_433 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(433), clk => clk, reset => reset); --
    end block;
    -- CP-element group 434:  transition  input  output  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	433 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	435 
    -- CP-element group 434:  members (6) 
      -- CP-element group 434: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1191_sample_completed_
      -- CP-element group 434: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1191_update_start_
      -- CP-element group 434: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1191_Sample/$exit
      -- CP-element group 434: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1191_Sample/ack
      -- CP-element group 434: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1191_Update/$entry
      -- CP-element group 434: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1191_Update/req
      -- 
    ack_2665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1191_inst_ack_0, ack => concat_CP_34_elements(434)); -- 
    req_2669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(434), ack => WPIPE_Concat_output_pipe_1191_inst_req_1); -- 
    -- CP-element group 435:  transition  input  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	434 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	436 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1191_update_completed_
      -- CP-element group 435: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1191_Update/$exit
      -- CP-element group 435: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/WPIPE_Concat_output_pipe_1191_Update/ack
      -- 
    ack_2670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1191_inst_ack_1, ack => concat_CP_34_elements(435)); -- 
    -- CP-element group 436:  branch  join  transition  place  output  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	391 
    -- CP-element group 436: 	435 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	437 
    -- CP-element group 436: 	438 
    -- CP-element group 436:  members (10) 
      -- CP-element group 436: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204__exit__
      -- CP-element group 436: 	 branch_block_stmt_23/if_stmt_1205__entry__
      -- CP-element group 436: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/$exit
      -- CP-element group 436: 	 branch_block_stmt_23/if_stmt_1205_dead_link/$entry
      -- CP-element group 436: 	 branch_block_stmt_23/if_stmt_1205_eval_test/$entry
      -- CP-element group 436: 	 branch_block_stmt_23/if_stmt_1205_eval_test/$exit
      -- CP-element group 436: 	 branch_block_stmt_23/if_stmt_1205_eval_test/branch_req
      -- CP-element group 436: 	 branch_block_stmt_23/R_exitcond1_1206_place
      -- CP-element group 436: 	 branch_block_stmt_23/if_stmt_1205_if_link/$entry
      -- CP-element group 436: 	 branch_block_stmt_23/if_stmt_1205_else_link/$entry
      -- 
    branch_req_2678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(436), ack => if_stmt_1205_branch_req_0); -- 
    concat_cp_element_group_436: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_436"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(391) & concat_CP_34_elements(435);
      gj_concat_cp_element_group_436 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(436), clk => clk, reset => reset); --
    end block;
    -- CP-element group 437:  merge  transition  place  input  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	436 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	459 
    -- CP-element group 437:  members (13) 
      -- CP-element group 437: 	 branch_block_stmt_23/merge_stmt_1211__exit__
      -- CP-element group 437: 	 branch_block_stmt_23/forx_xend456x_xloopexit_forx_xend456
      -- CP-element group 437: 	 branch_block_stmt_23/merge_stmt_1211_PhiReqMerge
      -- CP-element group 437: 	 branch_block_stmt_23/forx_xend456x_xloopexit_forx_xend456_PhiReq/$exit
      -- CP-element group 437: 	 branch_block_stmt_23/forx_xend456x_xloopexit_forx_xend456_PhiReq/$entry
      -- CP-element group 437: 	 branch_block_stmt_23/merge_stmt_1211_PhiAck/dummy
      -- CP-element group 437: 	 branch_block_stmt_23/merge_stmt_1211_PhiAck/$exit
      -- CP-element group 437: 	 branch_block_stmt_23/merge_stmt_1211_PhiAck/$entry
      -- CP-element group 437: 	 branch_block_stmt_23/forx_xbody383_forx_xend456x_xloopexit_PhiReq/$exit
      -- CP-element group 437: 	 branch_block_stmt_23/forx_xbody383_forx_xend456x_xloopexit_PhiReq/$entry
      -- CP-element group 437: 	 branch_block_stmt_23/if_stmt_1205_if_link/$exit
      -- CP-element group 437: 	 branch_block_stmt_23/if_stmt_1205_if_link/if_choice_transition
      -- CP-element group 437: 	 branch_block_stmt_23/forx_xbody383_forx_xend456x_xloopexit
      -- 
    if_choice_transition_2683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1205_branch_ack_1, ack => concat_CP_34_elements(437)); -- 
    -- CP-element group 438:  fork  transition  place  input  output  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	436 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	454 
    -- CP-element group 438: 	455 
    -- CP-element group 438:  members (12) 
      -- CP-element group 438: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/type_cast_1083/SplitProtocol/Sample/$entry
      -- CP-element group 438: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/$entry
      -- CP-element group 438: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/$entry
      -- CP-element group 438: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/type_cast_1083/SplitProtocol/$entry
      -- CP-element group 438: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/type_cast_1083/$entry
      -- CP-element group 438: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/$entry
      -- CP-element group 438: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/type_cast_1083/SplitProtocol/Sample/rr
      -- CP-element group 438: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/type_cast_1083/SplitProtocol/Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/type_cast_1083/SplitProtocol/Update/cr
      -- CP-element group 438: 	 branch_block_stmt_23/if_stmt_1205_else_link/$exit
      -- CP-element group 438: 	 branch_block_stmt_23/if_stmt_1205_else_link/else_choice_transition
      -- CP-element group 438: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383
      -- 
    else_choice_transition_2687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1205_branch_ack_0, ack => concat_CP_34_elements(438)); -- 
    rr_2885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(438), ack => type_cast_1083_inst_req_0); -- 
    cr_2890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(438), ack => type_cast_1083_inst_req_1); -- 
    -- CP-element group 439:  merge  branch  transition  place  output  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	133 
    -- CP-element group 439: 	88 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	89 
    -- CP-element group 439: 	90 
    -- CP-element group 439:  members (17) 
      -- CP-element group 439: 	 branch_block_stmt_23/merge_stmt_323__exit__
      -- CP-element group 439: 	 branch_block_stmt_23/assign_stmt_329__entry__
      -- CP-element group 439: 	 branch_block_stmt_23/assign_stmt_329__exit__
      -- CP-element group 439: 	 branch_block_stmt_23/if_stmt_330__entry__
      -- CP-element group 439: 	 branch_block_stmt_23/assign_stmt_329/$entry
      -- CP-element group 439: 	 branch_block_stmt_23/assign_stmt_329/$exit
      -- CP-element group 439: 	 branch_block_stmt_23/if_stmt_330_dead_link/$entry
      -- CP-element group 439: 	 branch_block_stmt_23/if_stmt_330_eval_test/$entry
      -- CP-element group 439: 	 branch_block_stmt_23/if_stmt_330_eval_test/$exit
      -- CP-element group 439: 	 branch_block_stmt_23/if_stmt_330_eval_test/branch_req
      -- CP-element group 439: 	 branch_block_stmt_23/R_cmp175463_331_place
      -- CP-element group 439: 	 branch_block_stmt_23/if_stmt_330_if_link/$entry
      -- CP-element group 439: 	 branch_block_stmt_23/if_stmt_330_else_link/$entry
      -- CP-element group 439: 	 branch_block_stmt_23/merge_stmt_323_PhiReqMerge
      -- CP-element group 439: 	 branch_block_stmt_23/merge_stmt_323_PhiAck/$entry
      -- CP-element group 439: 	 branch_block_stmt_23/merge_stmt_323_PhiAck/$exit
      -- CP-element group 439: 	 branch_block_stmt_23/merge_stmt_323_PhiAck/dummy
      -- 
    branch_req_698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(439), ack => if_stmt_330_branch_req_0); -- 
    concat_CP_34_elements(439) <= OrReduce(concat_CP_34_elements(133) & concat_CP_34_elements(88));
    -- CP-element group 440:  transition  output  delay-element  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	92 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	444 
    -- CP-element group 440:  members (5) 
      -- CP-element group 440: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/$exit
      -- CP-element group 440: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_374/$exit
      -- CP-element group 440: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/type_cast_378_konst_delay_trans
      -- CP-element group 440: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/$exit
      -- CP-element group 440: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_req
      -- 
    phi_stmt_374_req_2735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_374_req_2735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(440), ack => phi_stmt_374_req_0); -- 
    -- Element group concat_CP_34_elements(440) is a control-delay.
    cp_element_440_delay: control_delay_element  generic map(name => " 440_delay", delay_value => 1)  port map(req => concat_CP_34_elements(92), ack => concat_CP_34_elements(440), clk => clk, reset =>reset);
    -- CP-element group 441:  transition  input  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	134 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	443 
    -- CP-element group 441:  members (2) 
      -- CP-element group 441: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/type_cast_380/SplitProtocol/Sample/ra
      -- CP-element group 441: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/type_cast_380/SplitProtocol/Sample/$exit
      -- 
    ra_2755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_380_inst_ack_0, ack => concat_CP_34_elements(441)); -- 
    -- CP-element group 442:  transition  input  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	134 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	443 
    -- CP-element group 442:  members (2) 
      -- CP-element group 442: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/type_cast_380/SplitProtocol/Update/ca
      -- CP-element group 442: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/type_cast_380/SplitProtocol/Update/$exit
      -- 
    ca_2760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_380_inst_ack_1, ack => concat_CP_34_elements(442)); -- 
    -- CP-element group 443:  join  transition  output  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	441 
    -- CP-element group 443: 	442 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	444 
    -- CP-element group 443:  members (6) 
      -- CP-element group 443: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_req
      -- CP-element group 443: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 443: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/type_cast_380/SplitProtocol/$exit
      -- CP-element group 443: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/type_cast_380/$exit
      -- CP-element group 443: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/phi_stmt_374_sources/$exit
      -- CP-element group 443: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_374/$exit
      -- 
    phi_stmt_374_req_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_374_req_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(443), ack => phi_stmt_374_req_1); -- 
    concat_cp_element_group_443: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_443"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(441) & concat_CP_34_elements(442);
      gj_concat_cp_element_group_443 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(443), clk => clk, reset => reset); --
    end block;
    -- CP-element group 444:  merge  transition  place  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	440 
    -- CP-element group 444: 	443 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	445 
    -- CP-element group 444:  members (2) 
      -- CP-element group 444: 	 branch_block_stmt_23/merge_stmt_373_PhiAck/$entry
      -- CP-element group 444: 	 branch_block_stmt_23/merge_stmt_373_PhiReqMerge
      -- 
    concat_CP_34_elements(444) <= OrReduce(concat_CP_34_elements(440) & concat_CP_34_elements(443));
    -- CP-element group 445:  fork  transition  place  input  output  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	444 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	104 
    -- CP-element group 445: 	108 
    -- CP-element group 445: 	112 
    -- CP-element group 445: 	116 
    -- CP-element group 445: 	120 
    -- CP-element group 445: 	124 
    -- CP-element group 445: 	128 
    -- CP-element group 445: 	100 
    -- CP-element group 445: 	131 
    -- CP-element group 445: 	93 
    -- CP-element group 445: 	94 
    -- CP-element group 445: 	96 
    -- CP-element group 445: 	97 
    -- CP-element group 445:  members (56) 
      -- CP-element group 445: 	 branch_block_stmt_23/merge_stmt_373__exit__
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536__entry__
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_final_index_sum_regn_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_final_index_sum_regn_Update/req
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/addr_of_387_complete/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/addr_of_387_complete/req
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_390_sample_start_
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/addr_of_387_update_start_
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_index_resized_1
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_index_scaled_1
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_index_computed_1
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_index_resize_1/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_index_resize_1/$exit
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_index_resize_1/index_resize_req
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_index_resize_1/index_resize_ack
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_index_scale_1/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_index_scale_1/$exit
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_index_scale_1/scale_rename_req
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_index_scale_1/scale_rename_ack
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_final_index_sum_regn_update_start
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_final_index_sum_regn_Sample/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/array_obj_ref_386_final_index_sum_regn_Sample/req
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_390_Sample/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/RPIPE_Concat_input_pipe_390_Sample/rr
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_394_update_start_
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_394_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_394_Update/cr
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_407_update_start_
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_407_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_407_Update/cr
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_425_update_start_
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_425_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_425_Update/cr
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_443_update_start_
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_443_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_443_Update/cr
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_461_update_start_
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_461_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_461_Update/cr
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_479_update_start_
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_479_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_479_Update/cr
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_497_update_start_
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_497_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_497_Update/cr
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_515_update_start_
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_515_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/type_cast_515_Update/cr
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_update_start_
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Update/word_access_complete/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Update/word_access_complete/word_0/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/assign_stmt_388_to_assign_stmt_536/ptr_deref_523_Update/word_access_complete/word_0/cr
      -- CP-element group 445: 	 branch_block_stmt_23/merge_stmt_373_PhiAck/phi_stmt_374_ack
      -- CP-element group 445: 	 branch_block_stmt_23/merge_stmt_373_PhiAck/$exit
      -- 
    phi_stmt_374_ack_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_374_ack_0, ack => concat_CP_34_elements(445)); -- 
    req_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => array_obj_ref_386_index_offset_req_1); -- 
    req_774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => addr_of_387_final_reg_req_1); -- 
    req_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => array_obj_ref_386_index_offset_req_0); -- 
    rr_783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => RPIPE_Concat_input_pipe_390_inst_req_0); -- 
    cr_802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => type_cast_394_inst_req_1); -- 
    cr_830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => type_cast_407_inst_req_1); -- 
    cr_858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => type_cast_425_inst_req_1); -- 
    cr_886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => type_cast_443_inst_req_1); -- 
    cr_914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => type_cast_461_inst_req_1); -- 
    cr_942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => type_cast_479_inst_req_1); -- 
    cr_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => type_cast_497_inst_req_1); -- 
    cr_998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => type_cast_515_inst_req_1); -- 
    cr_1048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => ptr_deref_523_store_0_req_1); -- 
    -- CP-element group 446:  transition  output  delay-element  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	136 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	450 
    -- CP-element group 446:  members (5) 
      -- CP-element group 446: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/type_cast_585_konst_delay_trans
      -- CP-element group 446: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/$exit
      -- CP-element group 446: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_581/$exit
      -- CP-element group 446: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_req
      -- CP-element group 446: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/$exit
      -- 
    phi_stmt_581_req_2789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_581_req_2789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(446), ack => phi_stmt_581_req_0); -- 
    -- Element group concat_CP_34_elements(446) is a control-delay.
    cp_element_446_delay: control_delay_element  generic map(name => " 446_delay", delay_value => 1)  port map(req => concat_CP_34_elements(136), ack => concat_CP_34_elements(446), clk => clk, reset =>reset);
    -- CP-element group 447:  transition  input  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	178 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	449 
    -- CP-element group 447:  members (2) 
      -- CP-element group 447: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/type_cast_587/SplitProtocol/Sample/ra
      -- CP-element group 447: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/type_cast_587/SplitProtocol/Sample/$exit
      -- 
    ra_2809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_587_inst_ack_0, ack => concat_CP_34_elements(447)); -- 
    -- CP-element group 448:  transition  input  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	178 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (2) 
      -- CP-element group 448: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/type_cast_587/SplitProtocol/Update/ca
      -- CP-element group 448: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/type_cast_587/SplitProtocol/Update/$exit
      -- 
    ca_2814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_587_inst_ack_1, ack => concat_CP_34_elements(448)); -- 
    -- CP-element group 449:  join  transition  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	447 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	450 
    -- CP-element group 449:  members (6) 
      -- CP-element group 449: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/type_cast_587/SplitProtocol/$exit
      -- CP-element group 449: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_req
      -- CP-element group 449: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/$exit
      -- CP-element group 449: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/$exit
      -- CP-element group 449: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/$exit
      -- CP-element group 449: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_581/phi_stmt_581_sources/type_cast_587/$exit
      -- 
    phi_stmt_581_req_2815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_581_req_2815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(449), ack => phi_stmt_581_req_1); -- 
    concat_cp_element_group_449: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_449"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(447) & concat_CP_34_elements(448);
      gj_concat_cp_element_group_449 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 450:  merge  transition  place  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	446 
    -- CP-element group 450: 	449 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450:  members (2) 
      -- CP-element group 450: 	 branch_block_stmt_23/merge_stmt_580_PhiAck/$entry
      -- CP-element group 450: 	 branch_block_stmt_23/merge_stmt_580_PhiReqMerge
      -- 
    concat_CP_34_elements(450) <= OrReduce(concat_CP_34_elements(446) & concat_CP_34_elements(449));
    -- CP-element group 451:  fork  transition  place  input  output  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	175 
    -- CP-element group 451: 	160 
    -- CP-element group 451: 	172 
    -- CP-element group 451: 	168 
    -- CP-element group 451: 	137 
    -- CP-element group 451: 	138 
    -- CP-element group 451: 	140 
    -- CP-element group 451: 	141 
    -- CP-element group 451: 	144 
    -- CP-element group 451: 	148 
    -- CP-element group 451: 	152 
    -- CP-element group 451: 	156 
    -- CP-element group 451: 	164 
    -- CP-element group 451:  members (56) 
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_614_update_start_
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_686_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_614_Update/cr
      -- CP-element group 451: 	 branch_block_stmt_23/merge_stmt_580__exit__
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743__entry__
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_614_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_final_index_sum_regn_Sample/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_final_index_sum_regn_Update/req
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_final_index_sum_regn_update_start
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_final_index_sum_regn_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_704_update_start_
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_668_Update/cr
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_668_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/merge_stmt_580_PhiAck/phi_stmt_581_ack
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_686_update_start_
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_668_update_start_
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_update_start_
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_601_Update/cr
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_final_index_sum_regn_Sample/req
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_601_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_722_Update/cr
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_722_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/merge_stmt_580_PhiAck/$exit
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Update/word_access_complete/word_0/cr
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_601_update_start_
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Update/word_access_complete/word_0/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_632_Update/cr
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_632_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_722_update_start_
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_650_Update/cr
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_597_Sample/rr
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_650_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Update/word_access_complete/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_632_update_start_
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_597_Sample/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_index_scale_1/scale_rename_ack
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_index_scale_1/scale_rename_req
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_704_Update/cr
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/RPIPE_Concat_input_pipe_597_sample_start_
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_index_scale_1/$exit
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/addr_of_594_complete/req
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_704_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_index_scale_1/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_650_update_start_
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/addr_of_594_complete/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/ptr_deref_730_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/type_cast_686_Update/cr
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_index_resize_1/index_resize_ack
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_index_resize_1/index_resize_req
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_index_resize_1/$exit
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/$entry
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/addr_of_594_update_start_
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_index_resized_1
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_index_scaled_1
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_index_computed_1
      -- CP-element group 451: 	 branch_block_stmt_23/assign_stmt_595_to_assign_stmt_743/array_obj_ref_593_index_resize_1/$entry
      -- 
    phi_stmt_581_ack_2820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_581_ack_0, ack => concat_CP_34_elements(451)); -- 
    cr_1189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(451), ack => type_cast_614_inst_req_1); -- 
    req_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(451), ack => array_obj_ref_593_index_offset_req_1); -- 
    cr_1273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(451), ack => type_cast_668_inst_req_1); -- 
    cr_1161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(451), ack => type_cast_601_inst_req_1); -- 
    req_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(451), ack => array_obj_ref_593_index_offset_req_0); -- 
    cr_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(451), ack => type_cast_722_inst_req_1); -- 
    cr_1407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(451), ack => ptr_deref_730_store_0_req_1); -- 
    cr_1217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(451), ack => type_cast_632_inst_req_1); -- 
    cr_1245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(451), ack => type_cast_650_inst_req_1); -- 
    rr_1142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(451), ack => RPIPE_Concat_input_pipe_597_inst_req_0); -- 
    cr_1329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(451), ack => type_cast_704_inst_req_1); -- 
    req_1133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(451), ack => addr_of_594_final_reg_req_1); -- 
    cr_1301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(451), ack => type_cast_686_inst_req_1); -- 
    -- CP-element group 452:  merge  fork  transition  place  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	177 
    -- CP-element group 452: 	90 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	179 
    -- CP-element group 452: 	180 
    -- CP-element group 452:  members (13) 
      -- CP-element group 452: 	 branch_block_stmt_23/call_stmt_755/call_stmt_755_Update/ccr
      -- CP-element group 452: 	 branch_block_stmt_23/merge_stmt_752__exit__
      -- CP-element group 452: 	 branch_block_stmt_23/call_stmt_755__entry__
      -- CP-element group 452: 	 branch_block_stmt_23/call_stmt_755/call_stmt_755_Sample/crr
      -- CP-element group 452: 	 branch_block_stmt_23/call_stmt_755/call_stmt_755_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_23/call_stmt_755/call_stmt_755_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_23/call_stmt_755/call_stmt_755_update_start_
      -- CP-element group 452: 	 branch_block_stmt_23/call_stmt_755/call_stmt_755_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_23/call_stmt_755/$entry
      -- CP-element group 452: 	 branch_block_stmt_23/merge_stmt_752_PhiReqMerge
      -- CP-element group 452: 	 branch_block_stmt_23/merge_stmt_752_PhiAck/dummy
      -- CP-element group 452: 	 branch_block_stmt_23/merge_stmt_752_PhiAck/$exit
      -- CP-element group 452: 	 branch_block_stmt_23/merge_stmt_752_PhiAck/$entry
      -- 
    ccr_1443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(452), ack => call_stmt_755_call_req_1); -- 
    crr_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(452), ack => call_stmt_755_call_req_0); -- 
    concat_CP_34_elements(452) <= OrReduce(concat_CP_34_elements(177) & concat_CP_34_elements(90));
    -- CP-element group 453:  transition  output  delay-element  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	390 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	457 
    -- CP-element group 453:  members (5) 
      -- CP-element group 453: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_req
      -- CP-element group 453: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/type_cast_1081_konst_delay_trans
      -- CP-element group 453: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/$exit
      -- CP-element group 453: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/phi_stmt_1077/$exit
      -- CP-element group 453: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/$exit
      -- 
    phi_stmt_1077_req_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1077_req_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(453), ack => phi_stmt_1077_req_0); -- 
    -- Element group concat_CP_34_elements(453) is a control-delay.
    cp_element_453_delay: control_delay_element  generic map(name => " 453_delay", delay_value => 1)  port map(req => concat_CP_34_elements(390), ack => concat_CP_34_elements(453), clk => clk, reset =>reset);
    -- CP-element group 454:  transition  input  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	438 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	456 
    -- CP-element group 454:  members (2) 
      -- CP-element group 454: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/type_cast_1083/SplitProtocol/Sample/$exit
      -- CP-element group 454: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/type_cast_1083/SplitProtocol/Sample/ra
      -- 
    ra_2886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1083_inst_ack_0, ack => concat_CP_34_elements(454)); -- 
    -- CP-element group 455:  transition  input  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	438 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455:  members (2) 
      -- CP-element group 455: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/type_cast_1083/SplitProtocol/Update/$exit
      -- CP-element group 455: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/type_cast_1083/SplitProtocol/Update/ca
      -- 
    ca_2891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1083_inst_ack_1, ack => concat_CP_34_elements(455)); -- 
    -- CP-element group 456:  join  transition  output  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	454 
    -- CP-element group 456: 	455 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	457 
    -- CP-element group 456:  members (6) 
      -- CP-element group 456: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/$exit
      -- CP-element group 456: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/type_cast_1083/SplitProtocol/$exit
      -- CP-element group 456: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/$exit
      -- CP-element group 456: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_sources/type_cast_1083/$exit
      -- CP-element group 456: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/$exit
      -- CP-element group 456: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1077/phi_stmt_1077_req
      -- 
    phi_stmt_1077_req_2892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1077_req_2892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(456), ack => phi_stmt_1077_req_1); -- 
    concat_cp_element_group_456: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_456"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(454) & concat_CP_34_elements(455);
      gj_concat_cp_element_group_456 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(456), clk => clk, reset => reset); --
    end block;
    -- CP-element group 457:  merge  transition  place  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	453 
    -- CP-element group 457: 	456 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	458 
    -- CP-element group 457:  members (2) 
      -- CP-element group 457: 	 branch_block_stmt_23/merge_stmt_1076_PhiReqMerge
      -- CP-element group 457: 	 branch_block_stmt_23/merge_stmt_1076_PhiAck/$entry
      -- 
    concat_CP_34_elements(457) <= OrReduce(concat_CP_34_elements(453) & concat_CP_34_elements(456));
    -- CP-element group 458:  fork  transition  place  input  output  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	457 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	391 
    -- CP-element group 458: 	392 
    -- CP-element group 458: 	394 
    -- CP-element group 458: 	396 
    -- CP-element group 458: 	398 
    -- CP-element group 458: 	400 
    -- CP-element group 458: 	402 
    -- CP-element group 458: 	404 
    -- CP-element group 458: 	406 
    -- CP-element group 458: 	408 
    -- CP-element group 458: 	410 
    -- CP-element group 458: 	412 
    -- CP-element group 458:  members (53) 
      -- CP-element group 458: 	 branch_block_stmt_23/merge_stmt_1076__exit__
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204__entry__
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/addr_of_1090_update_start_
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_index_resized_1
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_index_scaled_1
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_index_computed_1
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_index_resize_1/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_index_resize_1/$exit
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_index_resize_1/index_resize_req
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_index_resize_1/index_resize_ack
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_index_scale_1/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_index_scale_1/$exit
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_index_scale_1/scale_rename_req
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_index_scale_1/scale_rename_ack
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_final_index_sum_regn_update_start
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_final_index_sum_regn_Sample/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_final_index_sum_regn_Sample/req
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_final_index_sum_regn_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/array_obj_ref_1089_final_index_sum_regn_Update/req
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/addr_of_1090_complete/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/addr_of_1090_complete/req
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_update_start_
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Update/word_access_complete/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Update/word_access_complete/word_0/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/ptr_deref_1094_Update/word_access_complete/word_0/cr
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1098_update_start_
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1098_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1098_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1108_update_start_
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1108_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1108_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1118_update_start_
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1118_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1118_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1128_update_start_
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1128_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1128_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1138_update_start_
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1138_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1138_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1148_update_start_
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1148_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1148_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1158_update_start_
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1158_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1158_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1168_update_start_
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1168_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/assign_stmt_1091_to_assign_stmt_1204/type_cast_1168_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_23/merge_stmt_1076_PhiAck/phi_stmt_1077_ack
      -- CP-element group 458: 	 branch_block_stmt_23/merge_stmt_1076_PhiAck/$exit
      -- 
    phi_stmt_1077_ack_2897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1077_ack_0, ack => concat_CP_34_elements(458)); -- 
    req_2375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(458), ack => array_obj_ref_1089_index_offset_req_0); -- 
    req_2380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(458), ack => array_obj_ref_1089_index_offset_req_1); -- 
    req_2395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(458), ack => addr_of_1090_final_reg_req_1); -- 
    cr_2440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(458), ack => ptr_deref_1094_load_0_req_1); -- 
    cr_2459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(458), ack => type_cast_1098_inst_req_1); -- 
    cr_2473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(458), ack => type_cast_1108_inst_req_1); -- 
    cr_2487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(458), ack => type_cast_1118_inst_req_1); -- 
    cr_2501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(458), ack => type_cast_1128_inst_req_1); -- 
    cr_2515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(458), ack => type_cast_1138_inst_req_1); -- 
    cr_2529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(458), ack => type_cast_1148_inst_req_1); -- 
    cr_2543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(458), ack => type_cast_1158_inst_req_1); -- 
    cr_2557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(458), ack => type_cast_1168_inst_req_1); -- 
    -- CP-element group 459:  merge  transition  place  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	388 
    -- CP-element group 459: 	437 
    -- CP-element group 459: successors 
    -- CP-element group 459:  members (16) 
      -- CP-element group 459: 	 $exit
      -- CP-element group 459: 	 branch_block_stmt_23/$exit
      -- CP-element group 459: 	 branch_block_stmt_23/branch_block_stmt_23__exit__
      -- CP-element group 459: 	 branch_block_stmt_23/merge_stmt_1213__exit__
      -- CP-element group 459: 	 branch_block_stmt_23/return__
      -- CP-element group 459: 	 branch_block_stmt_23/merge_stmt_1215__exit__
      -- CP-element group 459: 	 branch_block_stmt_23/merge_stmt_1213_PhiReqMerge
      -- CP-element group 459: 	 branch_block_stmt_23/merge_stmt_1215_PhiReqMerge
      -- CP-element group 459: 	 branch_block_stmt_23/merge_stmt_1215_PhiAck/dummy
      -- CP-element group 459: 	 branch_block_stmt_23/merge_stmt_1215_PhiAck/$exit
      -- CP-element group 459: 	 branch_block_stmt_23/merge_stmt_1215_PhiAck/$entry
      -- CP-element group 459: 	 branch_block_stmt_23/return___PhiReq/$exit
      -- CP-element group 459: 	 branch_block_stmt_23/return___PhiReq/$entry
      -- CP-element group 459: 	 branch_block_stmt_23/merge_stmt_1213_PhiAck/dummy
      -- CP-element group 459: 	 branch_block_stmt_23/merge_stmt_1213_PhiAck/$exit
      -- CP-element group 459: 	 branch_block_stmt_23/merge_stmt_1213_PhiAck/$entry
      -- 
    concat_CP_34_elements(459) <= OrReduce(concat_CP_34_elements(388) & concat_CP_34_elements(437));
    concat_do_while_stmt_784_terminator_2039: loop_terminator -- 
      generic map (name => " concat_do_while_stmt_784_terminator_2039", max_iterations_in_flight =>15) 
      port map(loop_body_exit => concat_CP_34_elements(185),loop_continue => concat_CP_34_elements(332),loop_terminate => concat_CP_34_elements(331),loop_back => concat_CP_34_elements(183),loop_exit => concat_CP_34_elements(182),clk => clk, reset => reset); -- 
    phi_stmt_786_phi_seq_1511_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(200);
      concat_CP_34_elements(203)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(203);
      concat_CP_34_elements(204)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(205);
      concat_CP_34_elements(201) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(198);
      concat_CP_34_elements(207)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(209);
      concat_CP_34_elements(208)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(210);
      concat_CP_34_elements(199) <= phi_mux_reqs(1);
      phi_stmt_786_phi_seq_1511 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_786_phi_seq_1511") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(190), 
          phi_sample_ack => concat_CP_34_elements(196), 
          phi_update_req => concat_CP_34_elements(192), 
          phi_update_ack => concat_CP_34_elements(197), 
          phi_mux_ack => concat_CP_34_elements(202), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_790_phi_seq_1555_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(219);
      concat_CP_34_elements(222)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(222);
      concat_CP_34_elements(223)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(224);
      concat_CP_34_elements(220) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(217);
      concat_CP_34_elements(226)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(228);
      concat_CP_34_elements(227)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(229);
      concat_CP_34_elements(218) <= phi_mux_reqs(1);
      phi_stmt_790_phi_seq_1555 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_790_phi_seq_1555") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(213), 
          phi_sample_ack => concat_CP_34_elements(214), 
          phi_update_req => concat_CP_34_elements(215), 
          phi_update_ack => concat_CP_34_elements(216), 
          phi_mux_ack => concat_CP_34_elements(221), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_794_phi_seq_1599_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(238);
      concat_CP_34_elements(241)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(241);
      concat_CP_34_elements(242)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(243);
      concat_CP_34_elements(239) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(236);
      concat_CP_34_elements(245)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(247);
      concat_CP_34_elements(246)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(248);
      concat_CP_34_elements(237) <= phi_mux_reqs(1);
      phi_stmt_794_phi_seq_1599 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_794_phi_seq_1599") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(232), 
          phi_sample_ack => concat_CP_34_elements(233), 
          phi_update_req => concat_CP_34_elements(234), 
          phi_update_ack => concat_CP_34_elements(235), 
          phi_mux_ack => concat_CP_34_elements(240), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_798_phi_seq_1643_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(257);
      concat_CP_34_elements(260)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(260);
      concat_CP_34_elements(261)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(262);
      concat_CP_34_elements(258) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(255);
      concat_CP_34_elements(264)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(266);
      concat_CP_34_elements(265)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(267);
      concat_CP_34_elements(256) <= phi_mux_reqs(1);
      phi_stmt_798_phi_seq_1643 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_798_phi_seq_1643") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(251), 
          phi_sample_ack => concat_CP_34_elements(252), 
          phi_update_req => concat_CP_34_elements(253), 
          phi_update_ack => concat_CP_34_elements(254), 
          phi_mux_ack => concat_CP_34_elements(259), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1463_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= concat_CP_34_elements(186);
        preds(1)  <= concat_CP_34_elements(187);
        entry_tmerge_1463 : transition_merge -- 
          generic map(name => " entry_tmerge_1463")
          port map (preds => preds, symbol_out => concat_CP_34_elements(188));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_876_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_883_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_892_wire : std_logic_vector(15 downto 0);
    signal MUX_859_wire : std_logic_vector(63 downto 0);
    signal NOT_u1_u1_907_wire : std_logic_vector(0 downto 0);
    signal R_indvar476_592_resized : std_logic_vector(13 downto 0);
    signal R_indvar476_592_scaled : std_logic_vector(13 downto 0);
    signal R_indvar489_385_resized : std_logic_vector(13 downto 0);
    signal R_indvar489_385_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1088_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1088_scaled : std_logic_vector(13 downto 0);
    signal SUB_u16_u16_853_853_delayed_1_0_865 : std_logic_vector(15 downto 0);
    signal SUB_u32_u32_891_891_delayed_1_0_904 : std_logic_vector(31 downto 0);
    signal ULT_u32_u1_910_wire : std_logic_vector(0 downto 0);
    signal add131_413 : std_logic_vector(63 downto 0);
    signal add137_431 : std_logic_vector(63 downto 0);
    signal add143_449 : std_logic_vector(63 downto 0);
    signal add149_467 : std_logic_vector(63 downto 0);
    signal add155_485 : std_logic_vector(63 downto 0);
    signal add161_503 : std_logic_vector(63 downto 0);
    signal add167_521 : std_logic_vector(63 downto 0);
    signal add187_620 : std_logic_vector(63 downto 0);
    signal add193_638 : std_logic_vector(63 downto 0);
    signal add199_656 : std_logic_vector(63 downto 0);
    signal add205_674 : std_logic_vector(63 downto 0);
    signal add211_692 : std_logic_vector(63 downto 0);
    signal add217_710 : std_logic_vector(63 downto 0);
    signal add223_728 : std_logic_vector(63 downto 0);
    signal add_inp1_790 : std_logic_vector(15 downto 0);
    signal add_inp1_init_770 : std_logic_vector(15 downto 0);
    signal add_inp2_794 : std_logic_vector(15 downto 0);
    signal add_inp2_init_774 : std_logic_vector(15 downto 0);
    signal add_out_786 : std_logic_vector(31 downto 0);
    signal add_out_init_766 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1089_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1089_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1089_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1089_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1089_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1089_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_386_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_386_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_386_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_386_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_386_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_386_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_593_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_593_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_593_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_593_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_593_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_593_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_813_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_813_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_813_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_813_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_813_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_813_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_829_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_829_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_829_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_829_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_829_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_829_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_845_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_845_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_845_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_845_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_845_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_845_root_address : std_logic_vector(13 downto 0);
    signal arrayidx227_595 : std_logic_vector(31 downto 0);
    signal arrayidx388_1091 : std_logic_vector(31 downto 0);
    signal arrayidx_388 : std_logic_vector(31 downto 0);
    signal call10_65 : std_logic_vector(7 downto 0);
    signal call124_391 : std_logic_vector(7 downto 0);
    signal call128_404 : std_logic_vector(7 downto 0);
    signal call134_422 : std_logic_vector(7 downto 0);
    signal call140_440 : std_logic_vector(7 downto 0);
    signal call146_458 : std_logic_vector(7 downto 0);
    signal call14_77 : std_logic_vector(7 downto 0);
    signal call152_476 : std_logic_vector(7 downto 0);
    signal call158_494 : std_logic_vector(7 downto 0);
    signal call164_512 : std_logic_vector(7 downto 0);
    signal call180_598 : std_logic_vector(7 downto 0);
    signal call184_611 : std_logic_vector(7 downto 0);
    signal call190_629 : std_logic_vector(7 downto 0);
    signal call196_647 : std_logic_vector(7 downto 0);
    signal call19_90 : std_logic_vector(7 downto 0);
    signal call202_665 : std_logic_vector(7 downto 0);
    signal call208_683 : std_logic_vector(7 downto 0);
    signal call214_701 : std_logic_vector(7 downto 0);
    signal call220_719 : std_logic_vector(7 downto 0);
    signal call233_755 : std_logic_vector(63 downto 0);
    signal call23_102 : std_logic_vector(7 downto 0);
    signal call28_115 : std_logic_vector(7 downto 0);
    signal call2_40 : std_logic_vector(7 downto 0);
    signal call310_917 : std_logic_vector(63 downto 0);
    signal call32_127 : std_logic_vector(7 downto 0);
    signal call37_140 : std_logic_vector(7 downto 0);
    signal call41_152 : std_logic_vector(7 downto 0);
    signal call46_165 : std_logic_vector(7 downto 0);
    signal call50_177 : std_logic_vector(7 downto 0);
    signal call55_191 : std_logic_vector(7 downto 0);
    signal call59_203 : std_logic_vector(7 downto 0);
    signal call5_52 : std_logic_vector(7 downto 0);
    signal call64_216 : std_logic_vector(7 downto 0);
    signal call68_228 : std_logic_vector(7 downto 0);
    signal call73_241 : std_logic_vector(7 downto 0);
    signal call_26 : std_logic_vector(7 downto 0);
    signal cmp175463_329 : std_logic_vector(0 downto 0);
    signal cmp381460_1038 : std_logic_vector(0 downto 0);
    signal cmp467_314 : std_logic_vector(0 downto 0);
    signal cmp_807 : std_logic_vector(0 downto 0);
    signal cmp_816_delayed_6_0_818 : std_logic_vector(0 downto 0);
    signal cmp_829_delayed_6_0_834 : std_logic_vector(0 downto 0);
    signal cmp_844_delayed_12_0_853 : std_logic_vector(0 downto 0);
    signal continue_flag_912 : std_logic_vector(0 downto 0);
    signal conv11_69 : std_logic_vector(15 downto 0);
    signal conv125_395 : std_logic_vector(63 downto 0);
    signal conv130_408 : std_logic_vector(63 downto 0);
    signal conv136_426 : std_logic_vector(63 downto 0);
    signal conv142_444 : std_logic_vector(63 downto 0);
    signal conv148_462 : std_logic_vector(63 downto 0);
    signal conv154_480 : std_logic_vector(63 downto 0);
    signal conv160_498 : std_logic_vector(63 downto 0);
    signal conv166_516 : std_logic_vector(63 downto 0);
    signal conv17_81 : std_logic_vector(15 downto 0);
    signal conv181_602 : std_logic_vector(63 downto 0);
    signal conv186_615 : std_logic_vector(63 downto 0);
    signal conv192_633 : std_logic_vector(63 downto 0);
    signal conv198_651 : std_logic_vector(63 downto 0);
    signal conv1_31 : std_logic_vector(15 downto 0);
    signal conv204_669 : std_logic_vector(63 downto 0);
    signal conv20_94 : std_logic_vector(15 downto 0);
    signal conv210_687 : std_logic_vector(63 downto 0);
    signal conv216_705 : std_logic_vector(63 downto 0);
    signal conv222_723 : std_logic_vector(63 downto 0);
    signal conv234_923 : std_logic_vector(63 downto 0);
    signal conv26_106 : std_logic_vector(15 downto 0);
    signal conv29_119 : std_logic_vector(15 downto 0);
    signal conv311_928 : std_logic_vector(63 downto 0);
    signal conv317_937 : std_logic_vector(7 downto 0);
    signal conv323_947 : std_logic_vector(7 downto 0);
    signal conv329_957 : std_logic_vector(7 downto 0);
    signal conv335_967 : std_logic_vector(7 downto 0);
    signal conv341_977 : std_logic_vector(7 downto 0);
    signal conv347_987 : std_logic_vector(7 downto 0);
    signal conv353_997 : std_logic_vector(7 downto 0);
    signal conv359_1007 : std_logic_vector(7 downto 0);
    signal conv35_131 : std_logic_vector(15 downto 0);
    signal conv38_144 : std_logic_vector(15 downto 0);
    signal conv393_1099 : std_logic_vector(7 downto 0);
    signal conv399_1109 : std_logic_vector(7 downto 0);
    signal conv3_44 : std_logic_vector(15 downto 0);
    signal conv405_1119 : std_logic_vector(7 downto 0);
    signal conv411_1129 : std_logic_vector(7 downto 0);
    signal conv417_1139 : std_logic_vector(7 downto 0);
    signal conv423_1149 : std_logic_vector(7 downto 0);
    signal conv429_1159 : std_logic_vector(7 downto 0);
    signal conv435_1169 : std_logic_vector(7 downto 0);
    signal conv44_156 : std_logic_vector(15 downto 0);
    signal conv47_169 : std_logic_vector(15 downto 0);
    signal conv53_182 : std_logic_vector(31 downto 0);
    signal conv56_195 : std_logic_vector(31 downto 0);
    signal conv62_207 : std_logic_vector(31 downto 0);
    signal conv65_220 : std_logic_vector(31 downto 0);
    signal conv71_232 : std_logic_vector(31 downto 0);
    signal conv74_245 : std_logic_vector(31 downto 0);
    signal conv8_56 : std_logic_vector(15 downto 0);
    signal count1_255 : std_logic_vector(15 downto 0);
    signal count2_273 : std_logic_vector(15 downto 0);
    signal count_inp1_798 : std_logic_vector(15 downto 0);
    signal count_inp1_init_778 : std_logic_vector(15 downto 0);
    signal exitcond1_1204 : std_logic_vector(0 downto 0);
    signal exitcond2_536 : std_logic_vector(0 downto 0);
    signal exitcond_743 : std_logic_vector(0 downto 0);
    signal i0_d0_49 : std_logic_vector(15 downto 0);
    signal i0_d1_74 : std_logic_vector(15 downto 0);
    signal i0_d2_99 : std_logic_vector(15 downto 0);
    signal i1_823 : std_logic_vector(63 downto 0);
    signal i1_d0_124 : std_logic_vector(15 downto 0);
    signal i1_d1_149 : std_logic_vector(15 downto 0);
    signal i1_d2_174 : std_logic_vector(15 downto 0);
    signal i2_839 : std_logic_vector(63 downto 0);
    signal iNsTr_19_358 : std_logic_vector(63 downto 0);
    signal iNsTr_32_565 : std_logic_vector(63 downto 0);
    signal iNsTr_79_1061 : std_logic_vector(63 downto 0);
    signal indvar476_581 : std_logic_vector(63 downto 0);
    signal indvar489_374 : std_logic_vector(63 downto 0);
    signal indvar_1077 : std_logic_vector(63 downto 0);
    signal indvarx_xnext477_738 : std_logic_vector(63 downto 0);
    signal indvarx_xnext490_531 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1199 : std_logic_vector(63 downto 0);
    signal inp0_d0_263 : std_logic_vector(31 downto 0);
    signal inp1_d0_281 : std_logic_vector(31 downto 0);
    signal inp1_mul_259 : std_logic_vector(31 downto 0);
    signal inp2_mul_277 : std_logic_vector(31 downto 0);
    signal input1_count_302 : std_logic_vector(15 downto 0);
    signal input1_size_268 : std_logic_vector(31 downto 0);
    signal input2_count_308 : std_logic_vector(15 downto 0);
    signal input2_size_286 : std_logic_vector(31 downto 0);
    signal iv1_815 : std_logic_vector(31 downto 0);
    signal iv2_831 : std_logic_vector(31 downto 0);
    signal konst_863_wire_constant : std_logic_vector(15 downto 0);
    signal konst_873_wire_constant : std_logic_vector(15 downto 0);
    signal konst_875_wire_constant : std_logic_vector(15 downto 0);
    signal konst_882_wire_constant : std_logic_vector(15 downto 0);
    signal konst_891_wire_constant : std_logic_vector(15 downto 0);
    signal konst_897_wire_constant : std_logic_vector(31 downto 0);
    signal konst_902_wire_constant : std_logic_vector(31 downto 0);
    signal mul100_291 : std_logic_vector(31 downto 0);
    signal my_flag_870 : std_logic_vector(0 downto 0);
    signal next_add_inp1_886 : std_logic_vector(15 downto 0);
    signal next_add_inp1_886_793_buffered : std_logic_vector(15 downto 0);
    signal next_add_inp2_894 : std_logic_vector(15 downto 0);
    signal next_add_inp2_894_797_buffered : std_logic_vector(15 downto 0);
    signal next_add_out_899 : std_logic_vector(31 downto 0);
    signal next_add_out_899_789_buffered : std_logic_vector(31 downto 0);
    signal next_count_inp1_878 : std_logic_vector(15 downto 0);
    signal next_count_inp1_878_801_buffered : std_logic_vector(15 downto 0);
    signal o0_200 : std_logic_vector(31 downto 0);
    signal o1_225 : std_logic_vector(31 downto 0);
    signal o2_250 : std_logic_vector(31 downto 0);
    signal out_concat_762 : std_logic_vector(31 downto 0);
    signal output_size_296 : std_logic_vector(31 downto 0);
    signal ov_842_delayed_7_0_850 : std_logic_vector(31 downto 0);
    signal ov_847 : std_logic_vector(31 downto 0);
    signal ptr_deref_1094_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1094_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1094_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1094_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1094_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_523_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_523_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_523_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_523_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_523_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_523_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_730_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_730_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_730_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_730_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_730_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_730_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_822_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_822_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_822_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_822_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_822_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_838_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_838_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_838_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_838_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_838_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_855_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_855_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_855_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_855_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_855_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_855_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl127_401 : std_logic_vector(63 downto 0);
    signal shl133_419 : std_logic_vector(63 downto 0);
    signal shl139_437 : std_logic_vector(63 downto 0);
    signal shl145_455 : std_logic_vector(63 downto 0);
    signal shl151_473 : std_logic_vector(63 downto 0);
    signal shl157_491 : std_logic_vector(63 downto 0);
    signal shl163_509 : std_logic_vector(63 downto 0);
    signal shl183_608 : std_logic_vector(63 downto 0);
    signal shl189_626 : std_logic_vector(63 downto 0);
    signal shl18_87 : std_logic_vector(15 downto 0);
    signal shl195_644 : std_logic_vector(63 downto 0);
    signal shl201_662 : std_logic_vector(63 downto 0);
    signal shl207_680 : std_logic_vector(63 downto 0);
    signal shl213_698 : std_logic_vector(63 downto 0);
    signal shl219_716 : std_logic_vector(63 downto 0);
    signal shl27_112 : std_logic_vector(15 downto 0);
    signal shl36_137 : std_logic_vector(15 downto 0);
    signal shl45_162 : std_logic_vector(15 downto 0);
    signal shl54_188 : std_logic_vector(31 downto 0);
    signal shl63_213 : std_logic_vector(31 downto 0);
    signal shl72_238 : std_logic_vector(31 downto 0);
    signal shl9_62 : std_logic_vector(15 downto 0);
    signal shl_37 : std_logic_vector(15 downto 0);
    signal shr320_943 : std_logic_vector(63 downto 0);
    signal shr326_953 : std_logic_vector(63 downto 0);
    signal shr332_963 : std_logic_vector(63 downto 0);
    signal shr338_973 : std_logic_vector(63 downto 0);
    signal shr344_983 : std_logic_vector(63 downto 0);
    signal shr350_993 : std_logic_vector(63 downto 0);
    signal shr356_1003 : std_logic_vector(63 downto 0);
    signal shr396_1105 : std_logic_vector(63 downto 0);
    signal shr402_1115 : std_logic_vector(63 downto 0);
    signal shr408_1125 : std_logic_vector(63 downto 0);
    signal shr414_1135 : std_logic_vector(63 downto 0);
    signal shr420_1145 : std_logic_vector(63 downto 0);
    signal shr426_1155 : std_logic_vector(63 downto 0);
    signal shr432_1165 : std_logic_vector(63 downto 0);
    signal sub_933 : std_logic_vector(63 downto 0);
    signal tmp389_1095 : std_logic_vector(63 downto 0);
    signal tmp471x_xop_1057 : std_logic_vector(31 downto 0);
    signal tmp472_1051 : std_logic_vector(0 downto 0);
    signal tmp475_1074 : std_logic_vector(63 downto 0);
    signal tmp482_549 : std_logic_vector(31 downto 0);
    signal tmp482x_xop_561 : std_logic_vector(31 downto 0);
    signal tmp483_555 : std_logic_vector(0 downto 0);
    signal tmp487_578 : std_logic_vector(63 downto 0);
    signal tmp495_342 : std_logic_vector(31 downto 0);
    signal tmp495x_xop_354 : std_logic_vector(31 downto 0);
    signal tmp496_348 : std_logic_vector(0 downto 0);
    signal tmp500_371 : std_logic_vector(63 downto 0);
    signal total_size_783 : std_logic_vector(15 downto 0);
    signal type_cast_1001_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1036_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1049_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1055_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1065_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1072_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1081_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1083_wire : std_logic_vector(63 downto 0);
    signal type_cast_1103_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_110_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1113_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1123_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1133_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1143_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1153_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1163_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1197_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_135_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_160_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_186_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_211_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_236_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_300_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_306_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_312_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_327_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_340_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_346_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_352_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_35_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_362_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_369_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_378_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_380_wire : std_logic_vector(63 downto 0);
    signal type_cast_399_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_417_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_435_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_453_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_471_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_489_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_507_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_529_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_547_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_553_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_559_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_569_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_576_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_585_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_587_wire : std_logic_vector(63 downto 0);
    signal type_cast_606_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_60_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_624_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_642_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_660_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_678_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_696_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_714_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_736_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_760_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_812_resized : std_logic_vector(13 downto 0);
    signal type_cast_812_scaled : std_logic_vector(13 downto 0);
    signal type_cast_812_wire : std_logic_vector(63 downto 0);
    signal type_cast_828_resized : std_logic_vector(13 downto 0);
    signal type_cast_828_scaled : std_logic_vector(13 downto 0);
    signal type_cast_828_wire : std_logic_vector(63 downto 0);
    signal type_cast_844_resized : std_logic_vector(13 downto 0);
    signal type_cast_844_scaled : std_logic_vector(13 downto 0);
    signal type_cast_844_wire : std_logic_vector(63 downto 0);
    signal type_cast_85_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_921_wire : std_logic_vector(63 downto 0);
    signal type_cast_926_wire : std_logic_vector(63 downto 0);
    signal type_cast_941_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_951_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_961_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_971_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_981_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_991_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop502_571 : std_logic_vector(63 downto 0);
    signal xx_xop503_364 : std_logic_vector(63 downto 0);
    signal xx_xop_1067 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    add_inp1_init_770 <= "0000000000000000";
    add_inp2_init_774 <= "0000000000000000";
    add_out_init_766 <= "00000000000000000000000000000000";
    array_obj_ref_1089_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1089_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1089_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1089_resized_base_address <= "00000000000000";
    array_obj_ref_386_constant_part_of_offset <= "00000000000000";
    array_obj_ref_386_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_386_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_386_resized_base_address <= "00000000000000";
    array_obj_ref_593_constant_part_of_offset <= "00000000000000";
    array_obj_ref_593_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_593_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_593_resized_base_address <= "00000000000000";
    array_obj_ref_813_constant_part_of_offset <= "00000000000000";
    array_obj_ref_813_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_813_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_813_resized_base_address <= "00000000000000";
    array_obj_ref_829_constant_part_of_offset <= "00000000000000";
    array_obj_ref_829_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_829_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_829_resized_base_address <= "00000000000000";
    array_obj_ref_845_constant_part_of_offset <= "00000000000000";
    array_obj_ref_845_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_845_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_845_resized_base_address <= "00000000000000";
    count_inp1_init_778 <= "0000000000000000";
    konst_863_wire_constant <= "0000000000000001";
    konst_873_wire_constant <= "0000000000000000";
    konst_875_wire_constant <= "0000000000000001";
    konst_882_wire_constant <= "0000000000000001";
    konst_891_wire_constant <= "0000000000000001";
    konst_897_wire_constant <= "00000000000000000000000000000001";
    konst_902_wire_constant <= "00000000000000000000000000000001";
    ptr_deref_1094_word_offset_0 <= "00000000000000";
    ptr_deref_523_word_offset_0 <= "00000000000000";
    ptr_deref_730_word_offset_0 <= "00000000000000";
    ptr_deref_822_word_offset_0 <= "00000000000000";
    ptr_deref_838_word_offset_0 <= "00000000000000";
    ptr_deref_855_word_offset_0 <= "00000000000000";
    type_cast_1001_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1036_wire_constant <= "00000000000000000000000000000111";
    type_cast_1049_wire_constant <= "00000000000000000000000000000001";
    type_cast_1055_wire_constant <= "11111111111111111111111111111111";
    type_cast_1065_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1072_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1081_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1103_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_110_wire_constant <= "0000000000001000";
    type_cast_1113_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1123_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1133_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1143_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1153_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1163_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1197_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_135_wire_constant <= "0000000000001000";
    type_cast_160_wire_constant <= "0000000000001000";
    type_cast_186_wire_constant <= "00000000000000000000000000001000";
    type_cast_211_wire_constant <= "00000000000000000000000000001000";
    type_cast_236_wire_constant <= "00000000000000000000000000001000";
    type_cast_300_wire_constant <= "0000000000000011";
    type_cast_306_wire_constant <= "0000000000000011";
    type_cast_312_wire_constant <= "00000000000000000000000000000111";
    type_cast_327_wire_constant <= "00000000000000000000000000000111";
    type_cast_340_wire_constant <= "00000000000000000000000000000011";
    type_cast_346_wire_constant <= "00000000000000000000000000000001";
    type_cast_352_wire_constant <= "11111111111111111111111111111111";
    type_cast_35_wire_constant <= "0000000000001000";
    type_cast_362_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_369_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_378_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_399_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_417_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_435_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_453_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_471_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_489_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_507_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_529_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_547_wire_constant <= "00000000000000000000000000000011";
    type_cast_553_wire_constant <= "00000000000000000000000000000001";
    type_cast_559_wire_constant <= "11111111111111111111111111111111";
    type_cast_569_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_576_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_585_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_606_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_60_wire_constant <= "0000000000001000";
    type_cast_624_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_642_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_660_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_678_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_696_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_714_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_736_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_760_wire_constant <= "00000000000000000000000000000011";
    type_cast_85_wire_constant <= "0000000000001000";
    type_cast_941_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_951_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_961_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_971_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_981_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_991_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    phi_stmt_1077: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1081_wire_constant & type_cast_1083_wire;
      req <= phi_stmt_1077_req_0 & phi_stmt_1077_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1077",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1077_ack_0,
          idata => idata,
          odata => indvar_1077,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1077
    phi_stmt_374: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_378_wire_constant & type_cast_380_wire;
      req <= phi_stmt_374_req_0 & phi_stmt_374_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_374",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_374_ack_0,
          idata => idata,
          odata => indvar489_374,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_374
    phi_stmt_581: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_585_wire_constant & type_cast_587_wire;
      req <= phi_stmt_581_req_0 & phi_stmt_581_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_581",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_581_ack_0,
          idata => idata,
          odata => indvar476_581,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_581
    phi_stmt_786: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_out_init_766 & next_add_out_899_789_buffered;
      req <= phi_stmt_786_req_0 & phi_stmt_786_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_786",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_786_ack_0,
          idata => idata,
          odata => add_out_786,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_786
    phi_stmt_790: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_inp1_init_770 & next_add_inp1_886_793_buffered;
      req <= phi_stmt_790_req_0 & phi_stmt_790_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_790",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_790_ack_0,
          idata => idata,
          odata => add_inp1_790,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_790
    phi_stmt_794: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_inp2_init_774 & next_add_inp2_894_797_buffered;
      req <= phi_stmt_794_req_0 & phi_stmt_794_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_794",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_794_ack_0,
          idata => idata,
          odata => add_inp2_794,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_794
    phi_stmt_798: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= count_inp1_init_778 & next_count_inp1_878_801_buffered;
      req <= phi_stmt_798_req_0 & phi_stmt_798_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_798",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_798_ack_0,
          idata => idata,
          odata => count_inp1_798,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_798
    -- flow-through select operator MUX_1073_inst
    tmp475_1074 <= xx_xop_1067 when (tmp472_1051(0) /=  '0') else type_cast_1072_wire_constant;
    -- flow-through select operator MUX_370_inst
    tmp500_371 <= xx_xop503_364 when (tmp496_348(0) /=  '0') else type_cast_369_wire_constant;
    -- flow-through select operator MUX_577_inst
    tmp487_578 <= xx_xop502_571 when (tmp483_555(0) /=  '0') else type_cast_576_wire_constant;
    MUX_859_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_859_inst_req_0;
      MUX_859_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_859_inst_req_1;
      MUX_859_inst_ack_1<= update_ack(0);
      MUX_859_inst: SelectSplitProtocol generic map(name => "MUX_859_inst", data_width => 64, buffering => 1, flow_through => false, full_rate => true) -- 
        port map( x => i1_823, y => i2_839, sel => cmp_844_delayed_12_0_853, z => MUX_859_wire, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_877_inst
    next_count_inp1_878 <= konst_873_wire_constant when (my_flag_870(0) /=  '0') else ADD_u16_u16_876_wire;
    -- flow-through select operator MUX_885_inst
    next_add_inp1_886 <= ADD_u16_u16_883_wire when (cmp_807(0) /=  '0') else add_inp1_790;
    -- flow-through select operator MUX_893_inst
    next_add_inp2_894 <= add_inp2_794 when (cmp_807(0) /=  '0') else ADD_u16_u16_892_wire;
    W_cmp_816_delayed_6_0_816_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_cmp_816_delayed_6_0_816_inst_req_0;
      W_cmp_816_delayed_6_0_816_inst_ack_0<= wack(0);
      rreq(0) <= W_cmp_816_delayed_6_0_816_inst_req_1;
      W_cmp_816_delayed_6_0_816_inst_ack_1<= rack(0);
      W_cmp_816_delayed_6_0_816_inst : InterlockBuffer generic map ( -- 
        name => "W_cmp_816_delayed_6_0_816_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp_807,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => cmp_816_delayed_6_0_818,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_cmp_829_delayed_6_0_832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_cmp_829_delayed_6_0_832_inst_req_0;
      W_cmp_829_delayed_6_0_832_inst_ack_0<= wack(0);
      rreq(0) <= W_cmp_829_delayed_6_0_832_inst_req_1;
      W_cmp_829_delayed_6_0_832_inst_ack_1<= rack(0);
      W_cmp_829_delayed_6_0_832_inst : InterlockBuffer generic map ( -- 
        name => "W_cmp_829_delayed_6_0_832_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp_807,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => cmp_829_delayed_6_0_834,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_cmp_844_delayed_12_0_851_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_cmp_844_delayed_12_0_851_inst_req_0;
      W_cmp_844_delayed_12_0_851_inst_ack_0<= wack(0);
      rreq(0) <= W_cmp_844_delayed_12_0_851_inst_req_1;
      W_cmp_844_delayed_12_0_851_inst_ack_1<= rack(0);
      W_cmp_844_delayed_12_0_851_inst : InterlockBuffer generic map ( -- 
        name => "W_cmp_844_delayed_12_0_851_inst",
        buffer_size => 12,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp_807,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => cmp_844_delayed_12_0_853,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ov_842_delayed_7_0_848_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ov_842_delayed_7_0_848_inst_req_0;
      W_ov_842_delayed_7_0_848_inst_ack_0<= wack(0);
      rreq(0) <= W_ov_842_delayed_7_0_848_inst_req_1;
      W_ov_842_delayed_7_0_848_inst_ack_1<= rack(0);
      W_ov_842_delayed_7_0_848_inst : InterlockBuffer generic map ( -- 
        name => "W_ov_842_delayed_7_0_848_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ov_847,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ov_842_delayed_7_0_850,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1090_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1090_final_reg_req_0;
      addr_of_1090_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1090_final_reg_req_1;
      addr_of_1090_final_reg_ack_1<= rack(0);
      addr_of_1090_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1090_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1089_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx388_1091,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_387_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_387_final_reg_req_0;
      addr_of_387_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_387_final_reg_req_1;
      addr_of_387_final_reg_ack_1<= rack(0);
      addr_of_387_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_387_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_386_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_388,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_594_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_594_final_reg_req_0;
      addr_of_594_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_594_final_reg_req_1;
      addr_of_594_final_reg_ack_1<= rack(0);
      addr_of_594_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_594_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_593_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx227_595,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_814_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_814_final_reg_req_0;
      addr_of_814_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_814_final_reg_req_1;
      addr_of_814_final_reg_ack_1<= rack(0);
      addr_of_814_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_814_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_813_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iv1_815,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_830_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_830_final_reg_req_0;
      addr_of_830_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_830_final_reg_req_1;
      addr_of_830_final_reg_ack_1<= rack(0);
      addr_of_830_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_830_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_829_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iv2_831,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_846_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_846_final_reg_req_0;
      addr_of_846_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_846_final_reg_req_1;
      addr_of_846_final_reg_ack_1<= rack(0);
      addr_of_846_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_846_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_845_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ov_847,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_inp1_886_793_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_inp1_886_793_buf_req_0;
      next_add_inp1_886_793_buf_ack_0<= wack(0);
      rreq(0) <= next_add_inp1_886_793_buf_req_1;
      next_add_inp1_886_793_buf_ack_1<= rack(0);
      next_add_inp1_886_793_buf : InterlockBuffer generic map ( -- 
        name => "next_add_inp1_886_793_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_inp1_886,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_inp1_886_793_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_inp2_894_797_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_inp2_894_797_buf_req_0;
      next_add_inp2_894_797_buf_ack_0<= wack(0);
      rreq(0) <= next_add_inp2_894_797_buf_req_1;
      next_add_inp2_894_797_buf_ack_1<= rack(0);
      next_add_inp2_894_797_buf : InterlockBuffer generic map ( -- 
        name => "next_add_inp2_894_797_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_inp2_894,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_inp2_894_797_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_out_899_789_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_out_899_789_buf_req_0;
      next_add_out_899_789_buf_ack_0<= wack(0);
      rreq(0) <= next_add_out_899_789_buf_req_1;
      next_add_out_899_789_buf_ack_1<= rack(0);
      next_add_out_899_789_buf : InterlockBuffer generic map ( -- 
        name => "next_add_out_899_789_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_out_899,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_out_899_789_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_count_inp1_878_801_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_inp1_878_801_buf_req_0;
      next_count_inp1_878_801_buf_ack_0<= wack(0);
      rreq(0) <= next_count_inp1_878_801_buf_req_1;
      next_count_inp1_878_801_buf_ack_1<= rack(0);
      next_count_inp1_878_801_buf : InterlockBuffer generic map ( -- 
        name => "next_count_inp1_878_801_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_inp1_878,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_inp1_878_801_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1006_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1006_inst_req_0;
      type_cast_1006_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1006_inst_req_1;
      type_cast_1006_inst_ack_1<= rack(0);
      type_cast_1006_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1006_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr356_1003,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv359_1007,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_105_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_105_inst_req_0;
      type_cast_105_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_105_inst_req_1;
      type_cast_105_inst_ack_1<= rack(0);
      type_cast_105_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_105_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_102,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_106,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1060_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1060_inst_req_0;
      type_cast_1060_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1060_inst_req_1;
      type_cast_1060_inst_ack_1<= rack(0);
      type_cast_1060_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1060_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp471x_xop_1057,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_79_1061,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1083_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1083_inst_req_0;
      type_cast_1083_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1083_inst_req_1;
      type_cast_1083_inst_ack_1<= rack(0);
      type_cast_1083_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1083_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1199,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1083_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1098_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1098_inst_req_0;
      type_cast_1098_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1098_inst_req_1;
      type_cast_1098_inst_ack_1<= rack(0);
      type_cast_1098_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1098_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp389_1095,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv393_1099,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1108_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1108_inst_req_0;
      type_cast_1108_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1108_inst_req_1;
      type_cast_1108_inst_ack_1<= rack(0);
      type_cast_1108_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1108_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr396_1105,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv399_1109,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1118_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1118_inst_req_0;
      type_cast_1118_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1118_inst_req_1;
      type_cast_1118_inst_ack_1<= rack(0);
      type_cast_1118_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1118_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr402_1115,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv405_1119,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1128_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1128_inst_req_0;
      type_cast_1128_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1128_inst_req_1;
      type_cast_1128_inst_ack_1<= rack(0);
      type_cast_1128_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1128_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr408_1125,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv411_1129,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1138_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1138_inst_req_0;
      type_cast_1138_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1138_inst_req_1;
      type_cast_1138_inst_ack_1<= rack(0);
      type_cast_1138_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1138_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr414_1135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv417_1139,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1148_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1148_inst_req_0;
      type_cast_1148_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1148_inst_req_1;
      type_cast_1148_inst_ack_1<= rack(0);
      type_cast_1148_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1148_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr420_1145,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv423_1149,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1158_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1158_inst_req_0;
      type_cast_1158_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1158_inst_req_1;
      type_cast_1158_inst_ack_1<= rack(0);
      type_cast_1158_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1158_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr426_1155,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv429_1159,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1168_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1168_inst_req_0;
      type_cast_1168_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1168_inst_req_1;
      type_cast_1168_inst_ack_1<= rack(0);
      type_cast_1168_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1168_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr432_1165,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv435_1169,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_118_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_118_inst_req_0;
      type_cast_118_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_118_inst_req_1;
      type_cast_118_inst_ack_1<= rack(0);
      type_cast_118_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_118_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_115,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_119,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_130_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_130_inst_req_0;
      type_cast_130_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_130_inst_req_1;
      type_cast_130_inst_ack_1<= rack(0);
      type_cast_130_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_130_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_127,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_131,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_143_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_143_inst_req_0;
      type_cast_143_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_143_inst_req_1;
      type_cast_143_inst_ack_1<= rack(0);
      type_cast_143_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_143_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_140,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_144,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_155_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_155_inst_req_0;
      type_cast_155_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_155_inst_req_1;
      type_cast_155_inst_ack_1<= rack(0);
      type_cast_155_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_155_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_152,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_156,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_168_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_168_inst_req_0;
      type_cast_168_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_168_inst_req_1;
      type_cast_168_inst_ack_1<= rack(0);
      type_cast_168_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_168_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_165,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_169,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_181_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_181_inst_req_0;
      type_cast_181_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_181_inst_req_1;
      type_cast_181_inst_ack_1<= rack(0);
      type_cast_181_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_181_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_177,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_182,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_194_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_194_inst_req_0;
      type_cast_194_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_194_inst_req_1;
      type_cast_194_inst_ack_1<= rack(0);
      type_cast_194_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_194_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_195,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_206_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_206_inst_req_0;
      type_cast_206_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_206_inst_req_1;
      type_cast_206_inst_ack_1<= rack(0);
      type_cast_206_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_206_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call59_203,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_207,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_219_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_219_inst_req_0;
      type_cast_219_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_219_inst_req_1;
      type_cast_219_inst_ack_1<= rack(0);
      type_cast_219_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_219_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call64_216,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_220,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_231_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_231_inst_req_0;
      type_cast_231_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_231_inst_req_1;
      type_cast_231_inst_ack_1<= rack(0);
      type_cast_231_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_231_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call68_228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_232,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_244_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_244_inst_req_0;
      type_cast_244_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_244_inst_req_1;
      type_cast_244_inst_ack_1<= rack(0);
      type_cast_244_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_244_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call73_241,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_245,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_258_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_258_inst_req_0;
      type_cast_258_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_258_inst_req_1;
      type_cast_258_inst_ack_1<= rack(0);
      type_cast_258_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_258_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count1_255,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inp1_mul_259,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_262_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_262_inst_req_0;
      type_cast_262_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_262_inst_req_1;
      type_cast_262_inst_ack_1<= rack(0);
      type_cast_262_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_262_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i0_d0_49,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inp0_d0_263,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_276_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_276_inst_req_0;
      type_cast_276_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_276_inst_req_1;
      type_cast_276_inst_ack_1<= rack(0);
      type_cast_276_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_276_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count2_273,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inp2_mul_277,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_280_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_280_inst_req_0;
      type_cast_280_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_280_inst_req_1;
      type_cast_280_inst_ack_1<= rack(0);
      type_cast_280_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_280_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1_d0_124,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inp1_d0_281,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_30_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_30_inst_req_0;
      type_cast_30_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_30_inst_req_1;
      type_cast_30_inst_ack_1<= rack(0);
      type_cast_30_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_30_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_26,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_31,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_357_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_357_inst_req_0;
      type_cast_357_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_357_inst_req_1;
      type_cast_357_inst_ack_1<= rack(0);
      type_cast_357_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_357_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp495x_xop_354,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_19_358,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_380_inst_req_0;
      type_cast_380_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_380_inst_req_1;
      type_cast_380_inst_ack_1<= rack(0);
      type_cast_380_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_380_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext490_531,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_380_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_394_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_394_inst_req_0;
      type_cast_394_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_394_inst_req_1;
      type_cast_394_inst_ack_1<= rack(0);
      type_cast_394_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_394_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_395,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_407_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_407_inst_req_0;
      type_cast_407_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_407_inst_req_1;
      type_cast_407_inst_ack_1<= rack(0);
      type_cast_407_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_407_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_404,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_408,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_425_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_425_inst_req_0;
      type_cast_425_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_425_inst_req_1;
      type_cast_425_inst_ack_1<= rack(0);
      type_cast_425_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_425_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call134_422,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv136_426,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_43_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_43_inst_req_0;
      type_cast_43_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_43_inst_req_1;
      type_cast_43_inst_ack_1<= rack(0);
      type_cast_43_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_43_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_40,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_44,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_443_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_443_inst_req_0;
      type_cast_443_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_443_inst_req_1;
      type_cast_443_inst_ack_1<= rack(0);
      type_cast_443_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_443_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call140_440,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv142_444,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_461_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_461_inst_req_0;
      type_cast_461_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_461_inst_req_1;
      type_cast_461_inst_ack_1<= rack(0);
      type_cast_461_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_461_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call146_458,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv148_462,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_479_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_479_inst_req_0;
      type_cast_479_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_479_inst_req_1;
      type_cast_479_inst_ack_1<= rack(0);
      type_cast_479_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_479_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call152_476,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv154_480,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_497_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_497_inst_req_0;
      type_cast_497_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_497_inst_req_1;
      type_cast_497_inst_ack_1<= rack(0);
      type_cast_497_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_497_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call158_494,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv160_498,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_515_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_515_inst_req_0;
      type_cast_515_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_515_inst_req_1;
      type_cast_515_inst_ack_1<= rack(0);
      type_cast_515_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_515_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv166_516,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_55_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_55_inst_req_0;
      type_cast_55_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_55_inst_req_1;
      type_cast_55_inst_ack_1<= rack(0);
      type_cast_55_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_55_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_52,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_56,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_564_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_564_inst_req_0;
      type_cast_564_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_564_inst_req_1;
      type_cast_564_inst_ack_1<= rack(0);
      type_cast_564_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_564_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp482x_xop_561,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_32_565,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_587_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_587_inst_req_0;
      type_cast_587_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_587_inst_req_1;
      type_cast_587_inst_ack_1<= rack(0);
      type_cast_587_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_587_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext477_738,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_587_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_601_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_601_inst_req_0;
      type_cast_601_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_601_inst_req_1;
      type_cast_601_inst_ack_1<= rack(0);
      type_cast_601_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_601_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call180_598,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv181_602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_614_inst_req_0;
      type_cast_614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_614_inst_req_1;
      type_cast_614_inst_ack_1<= rack(0);
      type_cast_614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call184_611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv186_615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_632_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_632_inst_req_0;
      type_cast_632_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_632_inst_req_1;
      type_cast_632_inst_ack_1<= rack(0);
      type_cast_632_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_632_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call190_629,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv192_633,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_650_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_650_inst_req_0;
      type_cast_650_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_650_inst_req_1;
      type_cast_650_inst_ack_1<= rack(0);
      type_cast_650_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_650_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call196_647,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv198_651,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_668_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_668_inst_req_0;
      type_cast_668_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_668_inst_req_1;
      type_cast_668_inst_ack_1<= rack(0);
      type_cast_668_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_668_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call202_665,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv204_669,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_686_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_686_inst_req_0;
      type_cast_686_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_686_inst_req_1;
      type_cast_686_inst_ack_1<= rack(0);
      type_cast_686_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_686_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call208_683,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv210_687,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_68_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_68_inst_req_0;
      type_cast_68_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_68_inst_req_1;
      type_cast_68_inst_ack_1<= rack(0);
      type_cast_68_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_68_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_65,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_69,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_704_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_704_inst_req_0;
      type_cast_704_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_704_inst_req_1;
      type_cast_704_inst_ack_1<= rack(0);
      type_cast_704_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_704_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call214_701,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv216_705,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_722_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_722_inst_req_0;
      type_cast_722_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_722_inst_req_1;
      type_cast_722_inst_ack_1<= rack(0);
      type_cast_722_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_722_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call220_719,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv222_723,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_80_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_80_inst_req_0;
      type_cast_80_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_80_inst_req_1;
      type_cast_80_inst_ack_1<= rack(0);
      type_cast_80_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_80_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_77,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_81,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_812_inst
    process(add_inp1_790) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := add_inp1_790(15 downto 0);
      type_cast_812_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_828_inst
    process(add_inp2_794) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := add_inp2_794(15 downto 0);
      type_cast_828_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_844_inst
    process(add_out_786) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_out_786(31 downto 0);
      type_cast_844_wire <= tmp_var; -- 
    end process;
    type_cast_922_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_922_inst_req_0;
      type_cast_922_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_922_inst_req_1;
      type_cast_922_inst_ack_1<= rack(0);
      type_cast_922_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_922_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_921_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv234_923,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_927_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_927_inst_req_0;
      type_cast_927_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_927_inst_req_1;
      type_cast_927_inst_ack_1<= rack(0);
      type_cast_927_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_927_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_926_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv311_928,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_936_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_936_inst_req_0;
      type_cast_936_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_936_inst_req_1;
      type_cast_936_inst_ack_1<= rack(0);
      type_cast_936_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_936_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_933,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv317_937,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_93_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_93_inst_req_0;
      type_cast_93_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_93_inst_req_1;
      type_cast_93_inst_ack_1<= rack(0);
      type_cast_93_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_93_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_90,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_94,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_946_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_946_inst_req_0;
      type_cast_946_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_946_inst_req_1;
      type_cast_946_inst_ack_1<= rack(0);
      type_cast_946_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_946_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr320_943,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv323_947,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_956_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_956_inst_req_0;
      type_cast_956_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_956_inst_req_1;
      type_cast_956_inst_ack_1<= rack(0);
      type_cast_956_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_956_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr326_953,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv329_957,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_966_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_966_inst_req_0;
      type_cast_966_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_966_inst_req_1;
      type_cast_966_inst_ack_1<= rack(0);
      type_cast_966_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_966_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr332_963,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv335_967,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_976_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_976_inst_req_0;
      type_cast_976_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_976_inst_req_1;
      type_cast_976_inst_ack_1<= rack(0);
      type_cast_976_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_976_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_973,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_977,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_986_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_986_inst_req_0;
      type_cast_986_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_986_inst_req_1;
      type_cast_986_inst_ack_1<= rack(0);
      type_cast_986_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_986_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr344_983,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv347_987,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_996_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_996_inst_req_0;
      type_cast_996_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_996_inst_req_1;
      type_cast_996_inst_ack_1<= rack(0);
      type_cast_996_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_996_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr350_993,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv353_997,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1089_index_1_rename
    process(R_indvar_1088_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1088_resized;
      ov(13 downto 0) := iv;
      R_indvar_1088_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1089_index_1_resize
    process(indvar_1077) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1077;
      ov := iv(13 downto 0);
      R_indvar_1088_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1089_root_address_inst
    process(array_obj_ref_1089_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1089_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1089_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_386_index_1_rename
    process(R_indvar489_385_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar489_385_resized;
      ov(13 downto 0) := iv;
      R_indvar489_385_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_386_index_1_resize
    process(indvar489_374) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar489_374;
      ov := iv(13 downto 0);
      R_indvar489_385_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_386_root_address_inst
    process(array_obj_ref_386_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_386_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_386_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_593_index_1_rename
    process(R_indvar476_592_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar476_592_resized;
      ov(13 downto 0) := iv;
      R_indvar476_592_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_593_index_1_resize
    process(indvar476_581) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar476_581;
      ov := iv(13 downto 0);
      R_indvar476_592_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_593_root_address_inst
    process(array_obj_ref_593_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_593_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_593_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_813_index_1_rename
    process(type_cast_812_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_812_resized;
      ov(13 downto 0) := iv;
      type_cast_812_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_813_index_1_resize
    process(type_cast_812_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_812_wire;
      ov := iv(13 downto 0);
      type_cast_812_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_813_root_address_inst
    process(array_obj_ref_813_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_813_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_813_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_829_index_1_rename
    process(type_cast_828_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_828_resized;
      ov(13 downto 0) := iv;
      type_cast_828_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_829_index_1_resize
    process(type_cast_828_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_828_wire;
      ov := iv(13 downto 0);
      type_cast_828_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_829_root_address_inst
    process(array_obj_ref_829_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_829_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_829_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_845_index_1_rename
    process(type_cast_844_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_844_resized;
      ov(13 downto 0) := iv;
      type_cast_844_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_845_index_1_resize
    process(type_cast_844_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_844_wire;
      ov := iv(13 downto 0);
      type_cast_844_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_845_root_address_inst
    process(array_obj_ref_845_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_845_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_845_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1094_addr_0
    process(ptr_deref_1094_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1094_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1094_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1094_base_resize
    process(arrayidx388_1091) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx388_1091;
      ov := iv(13 downto 0);
      ptr_deref_1094_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1094_gather_scatter
    process(ptr_deref_1094_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1094_data_0;
      ov(63 downto 0) := iv;
      tmp389_1095 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1094_root_address_inst
    process(ptr_deref_1094_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1094_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1094_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_523_addr_0
    process(ptr_deref_523_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_523_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_523_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_523_base_resize
    process(arrayidx_388) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_388;
      ov := iv(13 downto 0);
      ptr_deref_523_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_523_gather_scatter
    process(add167_521) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add167_521;
      ov(63 downto 0) := iv;
      ptr_deref_523_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_523_root_address_inst
    process(ptr_deref_523_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_523_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_523_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_730_addr_0
    process(ptr_deref_730_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_730_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_730_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_730_base_resize
    process(arrayidx227_595) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx227_595;
      ov := iv(13 downto 0);
      ptr_deref_730_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_730_gather_scatter
    process(add223_728) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add223_728;
      ov(63 downto 0) := iv;
      ptr_deref_730_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_730_root_address_inst
    process(ptr_deref_730_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_730_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_730_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_822_addr_0
    process(ptr_deref_822_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_822_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_822_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_822_base_resize
    process(iv1_815) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iv1_815;
      ov := iv(13 downto 0);
      ptr_deref_822_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_822_gather_scatter
    process(ptr_deref_822_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_822_data_0;
      ov(63 downto 0) := iv;
      i1_823 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_822_root_address_inst
    process(ptr_deref_822_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_822_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_822_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_838_addr_0
    process(ptr_deref_838_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_838_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_838_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_838_base_resize
    process(iv2_831) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iv2_831;
      ov := iv(13 downto 0);
      ptr_deref_838_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_838_gather_scatter
    process(ptr_deref_838_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_838_data_0;
      ov(63 downto 0) := iv;
      i2_839 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_838_root_address_inst
    process(ptr_deref_838_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_838_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_838_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_855_addr_0
    process(ptr_deref_855_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_855_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_855_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_855_base_resize
    process(ov_842_delayed_7_0_850) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ov_842_delayed_7_0_850;
      ov := iv(13 downto 0);
      ptr_deref_855_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_855_gather_scatter
    process(MUX_859_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := MUX_859_wire;
      ov(63 downto 0) := iv;
      ptr_deref_855_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_855_root_address_inst
    process(ptr_deref_855_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_855_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_855_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_784_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_912;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_784_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_784_branch_req_0,
          ack0 => do_while_stmt_784_branch_ack_0,
          ack1 => do_while_stmt_784_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1039_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp381460_1038;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1039_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1039_branch_req_0,
          ack0 => if_stmt_1039_branch_ack_0,
          ack1 => if_stmt_1039_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1205_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1204;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1205_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1205_branch_req_0,
          ack0 => if_stmt_1205_branch_ack_0,
          ack1 => if_stmt_1205_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_315_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp467_314;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_315_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_315_branch_req_0,
          ack0 => if_stmt_315_branch_ack_0,
          ack1 => if_stmt_315_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_330_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp175463_329;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_330_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_330_branch_req_0,
          ack0 => if_stmt_330_branch_ack_0,
          ack1 => if_stmt_330_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_537_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_536;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_537_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_537_branch_req_0,
          ack0 => if_stmt_537_branch_ack_0,
          ack1 => if_stmt_537_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_744_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_743;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_744_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_744_branch_req_0,
          ack0 => if_stmt_744_branch_ack_0,
          ack1 => if_stmt_744_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_782_inst
    process(input1_count_302, input2_count_308) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input1_count_302, input2_count_308, tmp_var);
      total_size_783 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_876_inst
    process(count_inp1_798) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(count_inp1_798, konst_875_wire_constant, tmp_var);
      ADD_u16_u16_876_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_883_inst
    process(add_inp1_790) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_inp1_790, konst_882_wire_constant, tmp_var);
      ADD_u16_u16_883_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_892_inst
    process(add_inp2_794) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_inp2_794, konst_891_wire_constant, tmp_var);
      ADD_u16_u16_892_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1056_inst
    process(out_concat_762) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(out_concat_762, type_cast_1055_wire_constant, tmp_var);
      tmp471x_xop_1057 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_353_inst
    process(tmp495_342) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp495_342, type_cast_352_wire_constant, tmp_var);
      tmp495x_xop_354 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_560_inst
    process(tmp482_549) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp482_549, type_cast_559_wire_constant, tmp_var);
      tmp482x_xop_561 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_898_inst
    process(add_out_786) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_out_786, konst_897_wire_constant, tmp_var);
      next_add_out_899 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1066_inst
    process(iNsTr_79_1061) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_79_1061, type_cast_1065_wire_constant, tmp_var);
      xx_xop_1067 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1198_inst
    process(indvar_1077) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1077, type_cast_1197_wire_constant, tmp_var);
      indvarx_xnext_1199 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_363_inst
    process(iNsTr_19_358) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_19_358, type_cast_362_wire_constant, tmp_var);
      xx_xop503_364 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_530_inst
    process(indvar489_374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar489_374, type_cast_529_wire_constant, tmp_var);
      indvarx_xnext490_531 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_570_inst
    process(iNsTr_32_565) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_32_565, type_cast_569_wire_constant, tmp_var);
      xx_xop502_571 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_737_inst
    process(indvar476_581) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar476_581, type_cast_736_wire_constant, tmp_var);
      indvarx_xnext477_738 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_869_inst
    process(count_inp1_798, SUB_u16_u16_853_853_delayed_1_0_865) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_inp1_798, SUB_u16_u16_853_853_delayed_1_0_865, tmp_var);
      my_flag_870 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1203_inst
    process(indvarx_xnext_1199, tmp475_1074) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1199, tmp475_1074, tmp_var);
      exitcond1_1204 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_535_inst
    process(indvarx_xnext490_531, tmp500_371) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext490_531, tmp500_371, tmp_var);
      exitcond2_536 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_742_inst
    process(indvarx_xnext477_738, tmp487_578) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext477_738, tmp487_578, tmp_var);
      exitcond_743 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_301_inst
    process(count1_255) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(count1_255, type_cast_300_wire_constant, tmp_var);
      input1_count_302 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_307_inst
    process(count2_273) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(count2_273, type_cast_306_wire_constant, tmp_var);
      input2_count_308 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_341_inst
    process(input1_size_268) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(input1_size_268, type_cast_340_wire_constant, tmp_var);
      tmp495_342 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_548_inst
    process(input2_size_286) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(input2_size_286, type_cast_547_wire_constant, tmp_var);
      tmp482_549 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_761_inst
    process(output_size_296) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(output_size_296, type_cast_760_wire_constant, tmp_var);
      out_concat_762 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1002_inst
    process(sub_933) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_933, type_cast_1001_wire_constant, tmp_var);
      shr356_1003 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1104_inst
    process(tmp389_1095) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1095, type_cast_1103_wire_constant, tmp_var);
      shr396_1105 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1114_inst
    process(tmp389_1095) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1095, type_cast_1113_wire_constant, tmp_var);
      shr402_1115 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1124_inst
    process(tmp389_1095) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1095, type_cast_1123_wire_constant, tmp_var);
      shr408_1125 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1134_inst
    process(tmp389_1095) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1095, type_cast_1133_wire_constant, tmp_var);
      shr414_1135 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1144_inst
    process(tmp389_1095) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1095, type_cast_1143_wire_constant, tmp_var);
      shr420_1145 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1154_inst
    process(tmp389_1095) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1095, type_cast_1153_wire_constant, tmp_var);
      shr426_1155 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1164_inst
    process(tmp389_1095) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1095, type_cast_1163_wire_constant, tmp_var);
      shr432_1165 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_942_inst
    process(sub_933) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_933, type_cast_941_wire_constant, tmp_var);
      shr320_943 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_952_inst
    process(sub_933) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_933, type_cast_951_wire_constant, tmp_var);
      shr326_953 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_962_inst
    process(sub_933) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_933, type_cast_961_wire_constant, tmp_var);
      shr332_963 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_972_inst
    process(sub_933) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_933, type_cast_971_wire_constant, tmp_var);
      shr338_973 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_982_inst
    process(sub_933) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_933, type_cast_981_wire_constant, tmp_var);
      shr344_983 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_992_inst
    process(sub_933) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_933, type_cast_991_wire_constant, tmp_var);
      shr350_993 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_254_inst
    process(i0_d1_74, i0_d2_99) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(i0_d1_74, i0_d2_99, tmp_var);
      count1_255 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_272_inst
    process(i1_d1_149, i1_d2_174) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(i1_d1_149, i1_d2_174, tmp_var);
      count2_273 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_267_inst
    process(inp1_mul_259, inp0_d0_263) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(inp1_mul_259, inp0_d0_263, tmp_var);
      input1_size_268 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_285_inst
    process(inp2_mul_277, inp1_d0_281) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(inp2_mul_277, inp1_d0_281, tmp_var);
      input2_size_286 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_290_inst
    process(o1_225, o2_250) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(o1_225, o2_250, tmp_var);
      mul100_291 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_295_inst
    process(mul100_291, o0_200) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul100_291, o0_200, tmp_var);
      output_size_296 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_907_inst
    process(my_flag_870) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", my_flag_870, tmp_var);
      NOT_u1_u1_907_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u16_u16_123_inst
    process(shl27_112, conv29_119) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_112, conv29_119, tmp_var);
      i1_d0_124 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_148_inst
    process(shl36_137, conv38_144) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_137, conv38_144, tmp_var);
      i1_d1_149 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_173_inst
    process(shl45_162, conv47_169) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_162, conv47_169, tmp_var);
      i1_d2_174 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_48_inst
    process(shl_37, conv3_44) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_37, conv3_44, tmp_var);
      i0_d0_49 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_73_inst
    process(shl9_62, conv11_69) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_62, conv11_69, tmp_var);
      i0_d1_74 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_98_inst
    process(shl18_87, conv20_94) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_87, conv20_94, tmp_var);
      i0_d2_99 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_911_inst
    process(NOT_u1_u1_907_wire, ULT_u32_u1_910_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_907_wire, ULT_u32_u1_910_wire, tmp_var);
      continue_flag_912 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_199_inst
    process(shl54_188, conv56_195) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_188, conv56_195, tmp_var);
      o0_200 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_224_inst
    process(shl63_213, conv65_220) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl63_213, conv65_220, tmp_var);
      o1_225 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_249_inst
    process(shl72_238, conv74_245) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl72_238, conv74_245, tmp_var);
      o2_250 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_412_inst
    process(shl127_401, conv130_408) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl127_401, conv130_408, tmp_var);
      add131_413 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_430_inst
    process(shl133_419, conv136_426) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl133_419, conv136_426, tmp_var);
      add137_431 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_448_inst
    process(shl139_437, conv142_444) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl139_437, conv142_444, tmp_var);
      add143_449 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_466_inst
    process(shl145_455, conv148_462) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl145_455, conv148_462, tmp_var);
      add149_467 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_484_inst
    process(shl151_473, conv154_480) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl151_473, conv154_480, tmp_var);
      add155_485 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_502_inst
    process(shl157_491, conv160_498) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl157_491, conv160_498, tmp_var);
      add161_503 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_520_inst
    process(shl163_509, conv166_516) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl163_509, conv166_516, tmp_var);
      add167_521 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_619_inst
    process(shl183_608, conv186_615) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl183_608, conv186_615, tmp_var);
      add187_620 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_637_inst
    process(shl189_626, conv192_633) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl189_626, conv192_633, tmp_var);
      add193_638 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_655_inst
    process(shl195_644, conv198_651) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl195_644, conv198_651, tmp_var);
      add199_656 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_673_inst
    process(shl201_662, conv204_669) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl201_662, conv204_669, tmp_var);
      add205_674 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_691_inst
    process(shl207_680, conv210_687) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl207_680, conv210_687, tmp_var);
      add211_692 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_709_inst
    process(shl213_698, conv216_705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl213_698, conv216_705, tmp_var);
      add217_710 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_727_inst
    process(shl219_716, conv222_723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl219_716, conv222_723, tmp_var);
      add223_728 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_111_inst
    process(conv26_106) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_106, type_cast_110_wire_constant, tmp_var);
      shl27_112 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_136_inst
    process(conv35_131) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_131, type_cast_135_wire_constant, tmp_var);
      shl36_137 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_161_inst
    process(conv44_156) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_156, type_cast_160_wire_constant, tmp_var);
      shl45_162 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_36_inst
    process(conv1_31) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_31, type_cast_35_wire_constant, tmp_var);
      shl_37 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_61_inst
    process(conv8_56) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_56, type_cast_60_wire_constant, tmp_var);
      shl9_62 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_86_inst
    process(conv17_81) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_81, type_cast_85_wire_constant, tmp_var);
      shl18_87 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_187_inst
    process(conv53_182) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_182, type_cast_186_wire_constant, tmp_var);
      shl54_188 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_212_inst
    process(conv62_207) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv62_207, type_cast_211_wire_constant, tmp_var);
      shl63_213 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_237_inst
    process(conv71_232) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv71_232, type_cast_236_wire_constant, tmp_var);
      shl72_238 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_400_inst
    process(conv125_395) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv125_395, type_cast_399_wire_constant, tmp_var);
      shl127_401 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_418_inst
    process(add131_413) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add131_413, type_cast_417_wire_constant, tmp_var);
      shl133_419 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_436_inst
    process(add137_431) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add137_431, type_cast_435_wire_constant, tmp_var);
      shl139_437 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_454_inst
    process(add143_449) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add143_449, type_cast_453_wire_constant, tmp_var);
      shl145_455 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_472_inst
    process(add149_467) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add149_467, type_cast_471_wire_constant, tmp_var);
      shl151_473 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_490_inst
    process(add155_485) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add155_485, type_cast_489_wire_constant, tmp_var);
      shl157_491 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_508_inst
    process(add161_503) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add161_503, type_cast_507_wire_constant, tmp_var);
      shl163_509 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_607_inst
    process(conv181_602) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv181_602, type_cast_606_wire_constant, tmp_var);
      shl183_608 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_625_inst
    process(add187_620) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add187_620, type_cast_624_wire_constant, tmp_var);
      shl189_626 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_643_inst
    process(add193_638) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add193_638, type_cast_642_wire_constant, tmp_var);
      shl195_644 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_661_inst
    process(add199_656) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add199_656, type_cast_660_wire_constant, tmp_var);
      shl201_662 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_679_inst
    process(add205_674) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add205_674, type_cast_678_wire_constant, tmp_var);
      shl207_680 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_697_inst
    process(add211_692) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add211_692, type_cast_696_wire_constant, tmp_var);
      shl213_698 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_715_inst
    process(add217_710) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add217_710, type_cast_714_wire_constant, tmp_var);
      shl219_716 <= tmp_var; --
    end process;
    -- shared split operator group (91) : SUB_u16_u16_864_inst 
    ApIntSub_group_91: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= total_size_783;
      SUB_u16_u16_853_853_delayed_1_0_865 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_864_inst_req_0;
      SUB_u16_u16_864_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_864_inst_req_1;
      SUB_u16_u16_864_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_91_gI: SplitGuardInterface generic map(name => "ApIntSub_group_91_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_91",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 91
    -- shared split operator group (92) : SUB_u32_u32_903_inst 
    ApIntSub_group_92: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= out_concat_762;
      SUB_u32_u32_891_891_delayed_1_0_904 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_903_inst_req_0;
      SUB_u32_u32_903_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_903_inst_req_1;
      SUB_u32_u32_903_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_92_gI: SplitGuardInterface generic map(name => "ApIntSub_group_92_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_92",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 92
    -- binary operator SUB_u64_u64_932_inst
    process(conv311_928, conv234_923) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv311_928, conv234_923, tmp_var);
      sub_933 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1037_inst
    process(output_size_296) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(output_size_296, type_cast_1036_wire_constant, tmp_var);
      cmp381460_1038 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1050_inst
    process(out_concat_762) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(out_concat_762, type_cast_1049_wire_constant, tmp_var);
      tmp472_1051 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_313_inst
    process(input1_size_268) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(input1_size_268, type_cast_312_wire_constant, tmp_var);
      cmp467_314 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_328_inst
    process(input2_size_286) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(input2_size_286, type_cast_327_wire_constant, tmp_var);
      cmp175463_329 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_347_inst
    process(tmp495_342) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp495_342, type_cast_346_wire_constant, tmp_var);
      tmp496_348 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_554_inst
    process(tmp482_549) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp482_549, type_cast_553_wire_constant, tmp_var);
      tmp483_555 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_806_inst
    process(count_inp1_798, input1_count_302) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(count_inp1_798, input1_count_302, tmp_var);
      cmp_807 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_910_inst
    process(add_out_786, SUB_u32_u32_891_891_delayed_1_0_904) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add_out_786, SUB_u32_u32_891_891_delayed_1_0_904, tmp_var);
      ULT_u32_u1_910_wire <= tmp_var; --
    end process;
    -- shared split operator group (102) : array_obj_ref_1089_index_offset 
    ApIntAdd_group_102: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1088_scaled;
      array_obj_ref_1089_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1089_index_offset_req_0;
      array_obj_ref_1089_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1089_index_offset_req_1;
      array_obj_ref_1089_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_102_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_102_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_102",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 102
    -- shared split operator group (103) : array_obj_ref_386_index_offset 
    ApIntAdd_group_103: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar489_385_scaled;
      array_obj_ref_386_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_386_index_offset_req_0;
      array_obj_ref_386_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_386_index_offset_req_1;
      array_obj_ref_386_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_103_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_103_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_103",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 103
    -- shared split operator group (104) : array_obj_ref_593_index_offset 
    ApIntAdd_group_104: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar476_592_scaled;
      array_obj_ref_593_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_593_index_offset_req_0;
      array_obj_ref_593_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_593_index_offset_req_1;
      array_obj_ref_593_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_104_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_104_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_104",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 104
    -- shared split operator group (105) : array_obj_ref_813_index_offset 
    ApIntAdd_group_105: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_812_scaled;
      array_obj_ref_813_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_813_index_offset_req_0;
      array_obj_ref_813_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_813_index_offset_req_1;
      array_obj_ref_813_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_105_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_105_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_105",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 105
    -- shared split operator group (106) : array_obj_ref_829_index_offset 
    ApIntAdd_group_106: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_828_scaled;
      array_obj_ref_829_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_829_index_offset_req_0;
      array_obj_ref_829_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_829_index_offset_req_1;
      array_obj_ref_829_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_106_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_106_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_106",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 106
    -- shared split operator group (107) : array_obj_ref_845_index_offset 
    ApIntAdd_group_107: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_844_scaled;
      array_obj_ref_845_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_845_index_offset_req_0;
      array_obj_ref_845_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_845_index_offset_req_1;
      array_obj_ref_845_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_107_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_107_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_107",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 107
    -- unary operator type_cast_921_inst
    process(call233_755) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call233_755, tmp_var);
      type_cast_921_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_926_inst
    process(call310_917) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call310_917, tmp_var);
      type_cast_926_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1094_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1094_load_0_req_0;
      ptr_deref_1094_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1094_load_0_req_1;
      ptr_deref_1094_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1094_word_address_0;
      ptr_deref_1094_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_822_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_822_load_0_req_0;
      ptr_deref_822_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_822_load_0_req_1;
      ptr_deref_822_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= cmp_816_delayed_6_0_818(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_822_word_address_0;
      ptr_deref_822_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_838_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_838_load_0_req_0;
      ptr_deref_838_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_838_load_0_req_1;
      ptr_deref_838_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not cmp_829_delayed_6_0_834(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_838_word_address_0;
      ptr_deref_838_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared store operator group (0) : ptr_deref_523_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_523_store_0_req_0;
      ptr_deref_523_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_523_store_0_req_1;
      ptr_deref_523_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_523_word_address_0;
      data_in <= ptr_deref_523_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_730_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_730_store_0_req_0;
      ptr_deref_730_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_730_store_0_req_1;
      ptr_deref_730_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_730_word_address_0;
      data_in <= ptr_deref_730_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_855_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 15);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_855_store_0_req_0;
      ptr_deref_855_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_855_store_0_req_1;
      ptr_deref_855_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_855_word_address_0;
      data_in <= ptr_deref_855_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Concat_input_pipe_439_inst RPIPE_Concat_input_pipe_664_inst RPIPE_Concat_input_pipe_421_inst RPIPE_Concat_input_pipe_390_inst RPIPE_Concat_input_pipe_457_inst RPIPE_Concat_input_pipe_240_inst RPIPE_Concat_input_pipe_646_inst RPIPE_Concat_input_pipe_682_inst RPIPE_Concat_input_pipe_610_inst RPIPE_Concat_input_pipe_215_inst RPIPE_Concat_input_pipe_718_inst RPIPE_Concat_input_pipe_700_inst RPIPE_Concat_input_pipe_403_inst RPIPE_Concat_input_pipe_227_inst RPIPE_Concat_input_pipe_597_inst RPIPE_Concat_input_pipe_628_inst RPIPE_Concat_input_pipe_493_inst RPIPE_Concat_input_pipe_475_inst RPIPE_Concat_input_pipe_511_inst RPIPE_Concat_input_pipe_25_inst RPIPE_Concat_input_pipe_39_inst RPIPE_Concat_input_pipe_51_inst RPIPE_Concat_input_pipe_64_inst RPIPE_Concat_input_pipe_76_inst RPIPE_Concat_input_pipe_89_inst RPIPE_Concat_input_pipe_101_inst RPIPE_Concat_input_pipe_114_inst RPIPE_Concat_input_pipe_126_inst RPIPE_Concat_input_pipe_139_inst RPIPE_Concat_input_pipe_151_inst RPIPE_Concat_input_pipe_164_inst RPIPE_Concat_input_pipe_176_inst RPIPE_Concat_input_pipe_190_inst RPIPE_Concat_input_pipe_202_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_Concat_input_pipe_439_inst_req_0;
      reqL_unguarded(32) <= RPIPE_Concat_input_pipe_664_inst_req_0;
      reqL_unguarded(31) <= RPIPE_Concat_input_pipe_421_inst_req_0;
      reqL_unguarded(30) <= RPIPE_Concat_input_pipe_390_inst_req_0;
      reqL_unguarded(29) <= RPIPE_Concat_input_pipe_457_inst_req_0;
      reqL_unguarded(28) <= RPIPE_Concat_input_pipe_240_inst_req_0;
      reqL_unguarded(27) <= RPIPE_Concat_input_pipe_646_inst_req_0;
      reqL_unguarded(26) <= RPIPE_Concat_input_pipe_682_inst_req_0;
      reqL_unguarded(25) <= RPIPE_Concat_input_pipe_610_inst_req_0;
      reqL_unguarded(24) <= RPIPE_Concat_input_pipe_215_inst_req_0;
      reqL_unguarded(23) <= RPIPE_Concat_input_pipe_718_inst_req_0;
      reqL_unguarded(22) <= RPIPE_Concat_input_pipe_700_inst_req_0;
      reqL_unguarded(21) <= RPIPE_Concat_input_pipe_403_inst_req_0;
      reqL_unguarded(20) <= RPIPE_Concat_input_pipe_227_inst_req_0;
      reqL_unguarded(19) <= RPIPE_Concat_input_pipe_597_inst_req_0;
      reqL_unguarded(18) <= RPIPE_Concat_input_pipe_628_inst_req_0;
      reqL_unguarded(17) <= RPIPE_Concat_input_pipe_493_inst_req_0;
      reqL_unguarded(16) <= RPIPE_Concat_input_pipe_475_inst_req_0;
      reqL_unguarded(15) <= RPIPE_Concat_input_pipe_511_inst_req_0;
      reqL_unguarded(14) <= RPIPE_Concat_input_pipe_25_inst_req_0;
      reqL_unguarded(13) <= RPIPE_Concat_input_pipe_39_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Concat_input_pipe_51_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Concat_input_pipe_64_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Concat_input_pipe_76_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Concat_input_pipe_89_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Concat_input_pipe_101_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Concat_input_pipe_114_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Concat_input_pipe_126_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Concat_input_pipe_139_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Concat_input_pipe_151_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Concat_input_pipe_164_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Concat_input_pipe_176_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Concat_input_pipe_190_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Concat_input_pipe_202_inst_req_0;
      RPIPE_Concat_input_pipe_439_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_Concat_input_pipe_664_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_Concat_input_pipe_421_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_Concat_input_pipe_390_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_Concat_input_pipe_457_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_Concat_input_pipe_240_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_Concat_input_pipe_646_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_Concat_input_pipe_682_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_Concat_input_pipe_610_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_Concat_input_pipe_215_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_Concat_input_pipe_718_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_Concat_input_pipe_700_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_Concat_input_pipe_403_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_Concat_input_pipe_227_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_Concat_input_pipe_597_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_Concat_input_pipe_628_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_Concat_input_pipe_493_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_Concat_input_pipe_475_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_Concat_input_pipe_511_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_Concat_input_pipe_25_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_Concat_input_pipe_39_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Concat_input_pipe_51_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Concat_input_pipe_64_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Concat_input_pipe_76_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Concat_input_pipe_89_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Concat_input_pipe_101_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Concat_input_pipe_114_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Concat_input_pipe_126_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Concat_input_pipe_139_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Concat_input_pipe_151_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Concat_input_pipe_164_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Concat_input_pipe_176_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Concat_input_pipe_190_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Concat_input_pipe_202_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_Concat_input_pipe_439_inst_req_1;
      reqR_unguarded(32) <= RPIPE_Concat_input_pipe_664_inst_req_1;
      reqR_unguarded(31) <= RPIPE_Concat_input_pipe_421_inst_req_1;
      reqR_unguarded(30) <= RPIPE_Concat_input_pipe_390_inst_req_1;
      reqR_unguarded(29) <= RPIPE_Concat_input_pipe_457_inst_req_1;
      reqR_unguarded(28) <= RPIPE_Concat_input_pipe_240_inst_req_1;
      reqR_unguarded(27) <= RPIPE_Concat_input_pipe_646_inst_req_1;
      reqR_unguarded(26) <= RPIPE_Concat_input_pipe_682_inst_req_1;
      reqR_unguarded(25) <= RPIPE_Concat_input_pipe_610_inst_req_1;
      reqR_unguarded(24) <= RPIPE_Concat_input_pipe_215_inst_req_1;
      reqR_unguarded(23) <= RPIPE_Concat_input_pipe_718_inst_req_1;
      reqR_unguarded(22) <= RPIPE_Concat_input_pipe_700_inst_req_1;
      reqR_unguarded(21) <= RPIPE_Concat_input_pipe_403_inst_req_1;
      reqR_unguarded(20) <= RPIPE_Concat_input_pipe_227_inst_req_1;
      reqR_unguarded(19) <= RPIPE_Concat_input_pipe_597_inst_req_1;
      reqR_unguarded(18) <= RPIPE_Concat_input_pipe_628_inst_req_1;
      reqR_unguarded(17) <= RPIPE_Concat_input_pipe_493_inst_req_1;
      reqR_unguarded(16) <= RPIPE_Concat_input_pipe_475_inst_req_1;
      reqR_unguarded(15) <= RPIPE_Concat_input_pipe_511_inst_req_1;
      reqR_unguarded(14) <= RPIPE_Concat_input_pipe_25_inst_req_1;
      reqR_unguarded(13) <= RPIPE_Concat_input_pipe_39_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Concat_input_pipe_51_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Concat_input_pipe_64_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Concat_input_pipe_76_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Concat_input_pipe_89_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Concat_input_pipe_101_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Concat_input_pipe_114_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Concat_input_pipe_126_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Concat_input_pipe_139_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Concat_input_pipe_151_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Concat_input_pipe_164_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Concat_input_pipe_176_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Concat_input_pipe_190_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Concat_input_pipe_202_inst_req_1;
      RPIPE_Concat_input_pipe_439_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_Concat_input_pipe_664_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_Concat_input_pipe_421_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_Concat_input_pipe_390_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_Concat_input_pipe_457_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_Concat_input_pipe_240_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_Concat_input_pipe_646_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_Concat_input_pipe_682_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_Concat_input_pipe_610_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_Concat_input_pipe_215_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_Concat_input_pipe_718_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_Concat_input_pipe_700_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_Concat_input_pipe_403_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_Concat_input_pipe_227_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_Concat_input_pipe_597_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_Concat_input_pipe_628_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_Concat_input_pipe_493_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_Concat_input_pipe_475_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_Concat_input_pipe_511_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_Concat_input_pipe_25_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_Concat_input_pipe_39_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Concat_input_pipe_51_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Concat_input_pipe_64_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Concat_input_pipe_76_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Concat_input_pipe_89_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Concat_input_pipe_101_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Concat_input_pipe_114_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Concat_input_pipe_126_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Concat_input_pipe_139_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Concat_input_pipe_151_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Concat_input_pipe_164_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Concat_input_pipe_176_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Concat_input_pipe_190_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Concat_input_pipe_202_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call140_440 <= data_out(271 downto 264);
      call202_665 <= data_out(263 downto 256);
      call134_422 <= data_out(255 downto 248);
      call124_391 <= data_out(247 downto 240);
      call146_458 <= data_out(239 downto 232);
      call73_241 <= data_out(231 downto 224);
      call196_647 <= data_out(223 downto 216);
      call208_683 <= data_out(215 downto 208);
      call184_611 <= data_out(207 downto 200);
      call64_216 <= data_out(199 downto 192);
      call220_719 <= data_out(191 downto 184);
      call214_701 <= data_out(183 downto 176);
      call128_404 <= data_out(175 downto 168);
      call68_228 <= data_out(167 downto 160);
      call180_598 <= data_out(159 downto 152);
      call190_629 <= data_out(151 downto 144);
      call158_494 <= data_out(143 downto 136);
      call152_476 <= data_out(135 downto 128);
      call164_512 <= data_out(127 downto 120);
      call_26 <= data_out(119 downto 112);
      call2_40 <= data_out(111 downto 104);
      call5_52 <= data_out(103 downto 96);
      call10_65 <= data_out(95 downto 88);
      call14_77 <= data_out(87 downto 80);
      call19_90 <= data_out(79 downto 72);
      call23_102 <= data_out(71 downto 64);
      call28_115 <= data_out(63 downto 56);
      call32_127 <= data_out(55 downto 48);
      call37_140 <= data_out(47 downto 40);
      call41_152 <= data_out(39 downto 32);
      call46_165 <= data_out(31 downto 24);
      call50_177 <= data_out(23 downto 16);
      call55_191 <= data_out(15 downto 8);
      call59_203 <= data_out(7 downto 0);
      Concat_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "Concat_input_pipe_read_0_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Concat_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "Concat_input_pipe_read_0", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Concat_input_pipe_pipe_read_req(0),
          oack => Concat_input_pipe_pipe_read_ack(0),
          odata => Concat_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Concat_output_pipe_1008_inst WPIPE_Concat_output_pipe_1011_inst WPIPE_Concat_output_pipe_1014_inst WPIPE_Concat_output_pipe_1017_inst WPIPE_Concat_output_pipe_1020_inst WPIPE_Concat_output_pipe_1023_inst WPIPE_Concat_output_pipe_1026_inst WPIPE_Concat_output_pipe_1029_inst WPIPE_Concat_output_pipe_1170_inst WPIPE_Concat_output_pipe_1173_inst WPIPE_Concat_output_pipe_1176_inst WPIPE_Concat_output_pipe_1179_inst WPIPE_Concat_output_pipe_1182_inst WPIPE_Concat_output_pipe_1185_inst WPIPE_Concat_output_pipe_1188_inst WPIPE_Concat_output_pipe_1191_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_Concat_output_pipe_1008_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_Concat_output_pipe_1011_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_Concat_output_pipe_1014_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Concat_output_pipe_1017_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Concat_output_pipe_1020_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Concat_output_pipe_1023_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Concat_output_pipe_1026_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Concat_output_pipe_1029_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Concat_output_pipe_1170_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Concat_output_pipe_1173_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Concat_output_pipe_1176_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Concat_output_pipe_1179_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Concat_output_pipe_1182_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Concat_output_pipe_1185_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Concat_output_pipe_1188_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Concat_output_pipe_1191_inst_req_0;
      WPIPE_Concat_output_pipe_1008_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_Concat_output_pipe_1011_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_Concat_output_pipe_1014_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Concat_output_pipe_1017_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Concat_output_pipe_1020_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Concat_output_pipe_1023_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Concat_output_pipe_1026_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Concat_output_pipe_1029_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Concat_output_pipe_1170_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Concat_output_pipe_1173_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Concat_output_pipe_1176_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Concat_output_pipe_1179_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Concat_output_pipe_1182_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Concat_output_pipe_1185_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Concat_output_pipe_1188_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Concat_output_pipe_1191_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_Concat_output_pipe_1008_inst_req_1;
      update_req_unguarded(14) <= WPIPE_Concat_output_pipe_1011_inst_req_1;
      update_req_unguarded(13) <= WPIPE_Concat_output_pipe_1014_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Concat_output_pipe_1017_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Concat_output_pipe_1020_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Concat_output_pipe_1023_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Concat_output_pipe_1026_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Concat_output_pipe_1029_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Concat_output_pipe_1170_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Concat_output_pipe_1173_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Concat_output_pipe_1176_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Concat_output_pipe_1179_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Concat_output_pipe_1182_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Concat_output_pipe_1185_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Concat_output_pipe_1188_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Concat_output_pipe_1191_inst_req_1;
      WPIPE_Concat_output_pipe_1008_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_Concat_output_pipe_1011_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_Concat_output_pipe_1014_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Concat_output_pipe_1017_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Concat_output_pipe_1020_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Concat_output_pipe_1023_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Concat_output_pipe_1026_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Concat_output_pipe_1029_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Concat_output_pipe_1170_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Concat_output_pipe_1173_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Concat_output_pipe_1176_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Concat_output_pipe_1179_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Concat_output_pipe_1182_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Concat_output_pipe_1185_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Concat_output_pipe_1188_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Concat_output_pipe_1191_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv359_1007 & conv353_997 & conv347_987 & conv341_977 & conv335_967 & conv329_957 & conv323_947 & conv317_937 & conv435_1169 & conv429_1159 & conv423_1149 & conv417_1139 & conv411_1129 & conv405_1119 & conv399_1109 & conv393_1099;
      Concat_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "Concat_output_pipe_write_0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Concat_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "Concat_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Concat_output_pipe_pipe_write_req(0),
          oack => Concat_output_pipe_pipe_write_ack(0),
          odata => Concat_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_755_call call_stmt_917_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_755_call_req_0;
      reqL_unguarded(0) <= call_stmt_917_call_req_0;
      call_stmt_755_call_ack_0 <= ackL_unguarded(1);
      call_stmt_917_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_755_call_req_1;
      reqR_unguarded(0) <= call_stmt_917_call_req_1;
      call_stmt_755_call_ack_1 <= ackR_unguarded(1);
      call_stmt_917_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call233_755 <= data_out(127 downto 64);
      call310_917 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end concat_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_14_inst_req_0 : boolean;
  signal WPIPE_timer_req_14_inst_ack_0 : boolean;
  signal WPIPE_timer_req_14_inst_req_1 : boolean;
  signal WPIPE_timer_req_14_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_19_inst_req_0 : boolean;
  signal RPIPE_timer_resp_19_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_19_inst_req_1 : boolean;
  signal RPIPE_timer_resp_19_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/$entry
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_sample_start_
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Sample/req
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_sample_start_
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Sample/rr
      -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => RPIPE_timer_resp_19_inst_req_0); -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => WPIPE_timer_req_14_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_sample_completed_
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_update_start_
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Sample/ack
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Update/$entry
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_14_inst_ack_0, ack => timer_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(1), ack => WPIPE_timer_req_14_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_update_completed_
      -- CP-element group 2: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Update/$exit
      -- CP-element group 2: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_14_inst_ack_1, ack => timer_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_update_start_
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_sample_completed_
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Sample/ra
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Update/$entry
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_19_inst_ack_0, ack => timer_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(3), ack => RPIPE_timer_resp_19_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_update_completed_
      -- CP-element group 4: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Update/$exit
      -- CP-element group 4: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_19_inst_ack_1, ack => timer_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_17_to_assign_stmt_20/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_0_elements(4) & timer_CP_0_elements(2);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_16_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_16_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_19_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_19_inst_req_0;
      RPIPE_timer_resp_19_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_19_inst_req_1;
      RPIPE_timer_resp_19_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_14_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_14_inst_req_0;
      WPIPE_timer_req_14_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_14_inst_req_1;
      WPIPE_timer_req_14_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_16_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_2932_start: Boolean;
  signal timerDaemon_CP_2932_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_resp_1240_inst_req_1 : boolean;
  signal WPIPE_timer_resp_1240_inst_ack_1 : boolean;
  signal phi_stmt_1225_ack_0 : boolean;
  signal do_while_stmt_1223_branch_req_0 : boolean;
  signal RPIPE_timer_req_1232_inst_req_0 : boolean;
  signal RPIPE_timer_req_1232_inst_ack_0 : boolean;
  signal nCOUNTER_1238_1229_buf_req_0 : boolean;
  signal nCOUNTER_1238_1229_buf_ack_0 : boolean;
  signal do_while_stmt_1223_branch_ack_0 : boolean;
  signal phi_stmt_1225_req_1 : boolean;
  signal phi_stmt_1225_req_0 : boolean;
  signal nCOUNTER_1238_1229_buf_req_1 : boolean;
  signal nCOUNTER_1238_1229_buf_ack_1 : boolean;
  signal RPIPE_timer_req_1232_inst_req_1 : boolean;
  signal do_while_stmt_1223_branch_ack_1 : boolean;
  signal WPIPE_timer_resp_1240_inst_req_0 : boolean;
  signal RPIPE_timer_req_1232_inst_ack_1 : boolean;
  signal WPIPE_timer_resp_1240_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_2932_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_2932_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_2932_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_2932_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_2932: Block -- control-path 
    signal timerDaemon_CP_2932_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_2932_elements(0) <= timerDaemon_CP_2932_start;
    timerDaemon_CP_2932_symbol <= timerDaemon_CP_2932_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1222/do_while_stmt_1223__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1222/branch_block_stmt_1222__entry__
      -- CP-element group 0: 	 branch_block_stmt_1222/$entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1222/do_while_stmt_1223__exit__
      -- CP-element group 1: 	 branch_block_stmt_1222/branch_block_stmt_1222__exit__
      -- CP-element group 1: 	 branch_block_stmt_1222/$exit
      -- 
    timerDaemon_CP_2932_elements(1) <= timerDaemon_CP_2932_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223__entry__
      -- CP-element group 2: 	 branch_block_stmt_1222/do_while_stmt_1223/$entry
      -- 
    timerDaemon_CP_2932_elements(2) <= timerDaemon_CP_2932_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223__exit__
      -- 
    -- Element group timerDaemon_CP_2932_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1222/do_while_stmt_1223/loop_back
      -- 
    -- Element group timerDaemon_CP_2932_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1222/do_while_stmt_1223/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1222/do_while_stmt_1223/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1222/do_while_stmt_1223/loop_taken/$entry
      -- 
    timerDaemon_CP_2932_elements(5) <= timerDaemon_CP_2932_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1222/do_while_stmt_1223/loop_body_done
      -- 
    timerDaemon_CP_2932_elements(6) <= timerDaemon_CP_2932_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_2932_elements(7) <= timerDaemon_CP_2932_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_2932_elements(8) <= timerDaemon_CP_2932_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	40 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1230_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/$entry
      -- 
    -- Element group timerDaemon_CP_2932_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	40 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/condition_evaluated
      -- 
    condition_evaluated_2956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2932_elements(10), ack => do_while_stmt_1223_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2932_elements(14) & timerDaemon_CP_2932_elements(40);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2932_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_2932_elements(9) & timerDaemon_CP_2932_elements(15) & timerDaemon_CP_2932_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2932_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1230_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2932_elements(17) & timerDaemon_CP_2932_elements(35);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2932_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2932_elements(16) & timerDaemon_CP_2932_elements(32);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2932_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2932_elements(18) & timerDaemon_CP_2932_elements(36);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2932_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2932_elements(9) & timerDaemon_CP_2932_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2932_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2932_elements(9) & timerDaemon_CP_2932_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2932_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_2932_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_2932_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_loopback_trigger
      -- 
    timerDaemon_CP_2932_elements(19) <= timerDaemon_CP_2932_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_loopback_sample_req_ps
      -- 
    phi_stmt_1225_loopback_sample_req_2971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1225_loopback_sample_req_2971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2932_elements(20), ack => phi_stmt_1225_req_1); -- 
    -- Element group timerDaemon_CP_2932_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_entry_trigger
      -- 
    timerDaemon_CP_2932_elements(21) <= timerDaemon_CP_2932_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_entry_sample_req_ps
      -- 
    phi_stmt_1225_entry_sample_req_2974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1225_entry_sample_req_2974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2932_elements(22), ack => phi_stmt_1225_req_0); -- 
    -- Element group timerDaemon_CP_2932_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1225_phi_mux_ack_ps
      -- 
    phi_stmt_1225_phi_mux_ack_2977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1225_ack_0, ack => timerDaemon_CP_2932_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/type_cast_1228_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/type_cast_1228_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/type_cast_1228_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/type_cast_1228_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_2932_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/type_cast_1228_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/type_cast_1228_update_start__ps
      -- 
    -- Element group timerDaemon_CP_2932_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/type_cast_1228_update_completed__ps
      -- 
    timerDaemon_CP_2932_elements(26) <= timerDaemon_CP_2932_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/type_cast_1228_update_completed_
      -- 
    -- Element group timerDaemon_CP_2932_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_2932_elements(25), ack => timerDaemon_CP_2932_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_Sample/req
      -- 
    req_2998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2932_elements(28), ack => nCOUNTER_1238_1229_buf_req_0); -- 
    -- Element group timerDaemon_CP_2932_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_Update/req
      -- 
    req_3003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2932_elements(29), ack => nCOUNTER_1238_1229_buf_req_1); -- 
    -- Element group timerDaemon_CP_2932_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_Sample/ack
      -- 
    ack_2999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1238_1229_buf_ack_0, ack => timerDaemon_CP_2932_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/R_nCOUNTER_1229_Update/ack
      -- 
    ack_3004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1238_1229_buf_ack_1, ack => timerDaemon_CP_2932_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1230_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2932_elements(9) & timerDaemon_CP_2932_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2932_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/RPIPE_timer_req_1232_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/RPIPE_timer_req_1232_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/RPIPE_timer_req_1232_sample_start_
      -- 
    rr_3017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2932_elements(33), ack => RPIPE_timer_req_1232_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2932_elements(11) & timerDaemon_CP_2932_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2932_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/RPIPE_timer_req_1232_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/RPIPE_timer_req_1232_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/RPIPE_timer_req_1232_update_start_
      -- 
    cr_3022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2932_elements(34), ack => RPIPE_timer_req_1232_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2932_elements(13) & timerDaemon_CP_2932_elements(35);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2932_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/RPIPE_timer_req_1232_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/RPIPE_timer_req_1232_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/RPIPE_timer_req_1232_sample_completed_
      -- 
    ra_3018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1232_inst_ack_0, ack => timerDaemon_CP_2932_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/RPIPE_timer_req_1232_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/phi_stmt_1230_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/RPIPE_timer_req_1232_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/RPIPE_timer_req_1232_update_completed_
      -- 
    ca_3023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1232_inst_ack_1, ack => timerDaemon_CP_2932_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	18 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/WPIPE_timer_resp_1240_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/WPIPE_timer_resp_1240_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/WPIPE_timer_resp_1240_sample_start_
      -- 
    req_3031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2932_elements(37), ack => WPIPE_timer_resp_1240_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_2932_elements(18) & timerDaemon_CP_2932_elements(36) & timerDaemon_CP_2932_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2932_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	16 
    -- CP-element group 38: 	32 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/WPIPE_timer_resp_1240_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/WPIPE_timer_resp_1240_Update/req
      -- CP-element group 38: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/WPIPE_timer_resp_1240_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/WPIPE_timer_resp_1240_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/WPIPE_timer_resp_1240_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/WPIPE_timer_resp_1240_sample_completed_
      -- 
    ack_3032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1240_inst_ack_0, ack => timerDaemon_CP_2932_elements(38)); -- 
    req_3036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2932_elements(38), ack => WPIPE_timer_resp_1240_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/WPIPE_timer_resp_1240_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/WPIPE_timer_resp_1240_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/WPIPE_timer_resp_1240_Update/$exit
      -- 
    ack_3037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1240_inst_ack_1, ack => timerDaemon_CP_2932_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_2932_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_2932_elements(9), ack => timerDaemon_CP_2932_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	12 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1222/do_while_stmt_1223/do_while_stmt_1223_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2932_elements(12) & timerDaemon_CP_2932_elements(39);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2932_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1222/do_while_stmt_1223/loop_exit/$exit
      -- CP-element group 42: 	 branch_block_stmt_1222/do_while_stmt_1223/loop_exit/ack
      -- 
    ack_3042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1223_branch_ack_0, ack => timerDaemon_CP_2932_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1222/do_while_stmt_1223/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_1222/do_while_stmt_1223/loop_taken/ack
      -- 
    ack_3046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1223_branch_ack_1, ack => timerDaemon_CP_2932_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1222/do_while_stmt_1223/$exit
      -- 
    timerDaemon_CP_2932_elements(44) <= timerDaemon_CP_2932_elements(3);
    timerDaemon_do_while_stmt_1223_terminator_3047: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_1223_terminator_3047", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_2932_elements(6),loop_continue => timerDaemon_CP_2932_elements(43),loop_terminate => timerDaemon_CP_2932_elements(42),loop_back => timerDaemon_CP_2932_elements(4),loop_exit => timerDaemon_CP_2932_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1225_phi_seq_3005_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_2932_elements(21);
      timerDaemon_CP_2932_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_2932_elements(24);
      timerDaemon_CP_2932_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_2932_elements(26);
      timerDaemon_CP_2932_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_2932_elements(19);
      timerDaemon_CP_2932_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_2932_elements(30);
      timerDaemon_CP_2932_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_2932_elements(31);
      timerDaemon_CP_2932_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1225_phi_seq_3005 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1225_phi_seq_3005") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_2932_elements(11), 
          phi_sample_ack => timerDaemon_CP_2932_elements(17), 
          phi_update_req => timerDaemon_CP_2932_elements(13), 
          phi_update_ack => timerDaemon_CP_2932_elements(18), 
          phi_mux_ack => timerDaemon_CP_2932_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2957_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_2932_elements(7);
        preds(1)  <= timerDaemon_CP_2932_elements(8);
        entry_tmerge_2957 : transition_merge -- 
          generic map(name => " entry_tmerge_2957")
          port map (preds => preds, symbol_out => timerDaemon_CP_2932_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_1225 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_1232_wire : std_logic_vector(0 downto 0);
    signal konst_1236_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1244_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_1238 : std_logic_vector(63 downto 0);
    signal nCOUNTER_1238_1229_buffered : std_logic_vector(63 downto 0);
    signal req_1230 : std_logic_vector(0 downto 0);
    signal type_cast_1228_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_1236_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_1244_wire_constant <= "1";
    type_cast_1228_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1225: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1228_wire_constant & nCOUNTER_1238_1229_buffered;
      req <= phi_stmt_1225_req_0 & phi_stmt_1225_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1225",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1225_ack_0,
          idata => idata,
          odata => COUNTER_1225,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1225
    nCOUNTER_1238_1229_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_1238_1229_buf_req_0;
      nCOUNTER_1238_1229_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_1238_1229_buf_req_1;
      nCOUNTER_1238_1229_buf_ack_1<= rack(0);
      nCOUNTER_1238_1229_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_1238_1229_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_1238,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_1238_1229_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1230
    process(RPIPE_timer_req_1232_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_1232_wire(0 downto 0);
      req_1230 <= tmp_var; -- 
    end process;
    do_while_stmt_1223_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1244_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1223_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1223_branch_req_0,
          ack0 => do_while_stmt_1223_branch_ack_0,
          ack1 => do_while_stmt_1223_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_1237_inst
    process(COUNTER_1225) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_1225, konst_1236_wire_constant, tmp_var);
      nCOUNTER_1238 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_1232_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_1232_inst_req_0;
      RPIPE_timer_req_1232_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_1232_inst_req_1;
      RPIPE_timer_req_1232_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_1232_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_1240_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_1240_inst_req_0;
      WPIPE_timer_resp_1240_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_1240_inst_req_1;
      WPIPE_timer_resp_1240_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_1230(0);
      data_in <= COUNTER_1225;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    Concat_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    Concat_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    Concat_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    Concat_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module concat
  component concat is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      Concat_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      Concat_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Concat_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Concat_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      Concat_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Concat_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module concat
  signal concat_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal concat_tag_out   : std_logic_vector(1 downto 0);
  signal concat_start_req : std_logic;
  signal concat_start_ack : std_logic;
  signal concat_fin_req   : std_logic;
  signal concat_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for read from pipe Concat_input_pipe
  signal Concat_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal Concat_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal Concat_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Concat_output_pipe
  signal Concat_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal Concat_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal Concat_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module concat
  concat_instance:concat-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => concat_start_req,
      start_ack => concat_start_ack,
      fin_req => concat_fin_req,
      fin_ack => concat_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(17 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(17 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(17 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(17 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      Concat_input_pipe_pipe_read_req => Concat_input_pipe_pipe_read_req(0 downto 0),
      Concat_input_pipe_pipe_read_ack => Concat_input_pipe_pipe_read_ack(0 downto 0),
      Concat_input_pipe_pipe_read_data => Concat_input_pipe_pipe_read_data(7 downto 0),
      Concat_output_pipe_pipe_write_req => Concat_output_pipe_pipe_write_req(0 downto 0),
      Concat_output_pipe_pipe_write_ack => Concat_output_pipe_pipe_write_ack(0 downto 0),
      Concat_output_pipe_pipe_write_data => Concat_output_pipe_pipe_write_data(7 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => concat_tag_in,
      tag_out => concat_tag_out-- 
    ); -- 
  -- module will be run forever 
  concat_tag_in <= (others => '0');
  concat_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => concat_start_req, start_ack => concat_start_ack,  fin_req => concat_fin_req,  fin_ack => concat_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  Concat_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Concat_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => Concat_input_pipe_pipe_read_req,
      read_ack => Concat_input_pipe_pipe_read_ack,
      read_data => Concat_input_pipe_pipe_read_data,
      write_req => Concat_input_pipe_pipe_write_req,
      write_ack => Concat_input_pipe_pipe_write_ack,
      write_data => Concat_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Concat_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Concat_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => Concat_output_pipe_pipe_read_req,
      read_ack => Concat_output_pipe_pipe_read_ack,
      read_data => Concat_output_pipe_pipe_read_data,
      write_req => Concat_output_pipe_pipe_write_req,
      write_ack => Concat_output_pipe_pipe_write_ack,
      write_data => Concat_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
